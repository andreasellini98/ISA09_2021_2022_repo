LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;

ENTITY dadda IS
	GENERIC( NB: integer:= 32);
	PORT(
		a		: IN  std_logic_vector(NB-1 downto 0);
		b		: IN  std_logic_vector(NB-1 downto 0);
		prod	: OUT std_logic_vector(2*NB-1 downto 0)
	);
END ENTITY;

ARCHITECTURE struct OF dadda IS

COMPONENT MBE IS
	GENERIC ( NB : NATURAL := 32 );
	PORT( 
		a	: IN  std_logic_vector(NB-1 downto 0);
		b  	: IN  std_logic_vector(2 downto 0);
		p : OUT std_logic_vector(NB downto 0)
   );
END COMPONENT;

COMPONENT Half_Adder IS
PORT (
	a : IN STD_LOGIC;
	b : IN STD_LOGIC;
	s : OUT STD_LOGIC;
	cout : OUT STD_LOGIC
);
END COMPONENT;

COMPONENT Full_Adder IS
PORT (
	a 		: IN STD_LOGIC;
	b 		: IN STD_LOGIC;
	cin 	: IN STD_LOGIC;
	s 		: OUT STD_LOGIC;
	cout	: OUT STD_LOGIC
);
END COMPONENT;

COMPONENT ks_adder IS
	GENERIC( N: integer:= 64);
	PORT(
		a		: IN  std_logic_vector(N-1 downto 0);
		b		: IN  std_logic_vector(N-1 downto 0);
		sum		: OUT std_logic_vector(N-1 downto 0)
	);
END COMPONENT;


TYPE pptype IS ARRAY(0 to NB/2) OF std_logic_vector(NB DOWNTO 0);

TYPE p_layer_0 IS ARRAY(0 to 1) OF STD_LOGIC_VECTOR(2*NB DOWNTO 0); 
TYPE p_layer_1 IS ARRAY(0 to 2) OF STD_LOGIC_VECTOR(2*NB-1 DOWNTO 0); 
TYPE p_layer_2 IS ARRAY(0 to 3) OF STD_LOGIC_VECTOR(2*NB-1 DOWNTO 0); 
TYPE p_layer_3 IS ARRAY(0 to 5) OF STD_LOGIC_VECTOR(2*NB-1 DOWNTO 0); 
TYPE p_layer_4 IS ARRAY(0 to 8) OF STD_LOGIC_VECTOR(2*NB-1 DOWNTO 0); 
TYPE p_layer_5 IS ARRAY(0 to 12) OF STD_LOGIC_VECTOR(2*NB-1 DOWNTO 0); 
TYPE p_layer_6 IS ARRAY(0 to 16) OF STD_LOGIC_VECTOR(2*NB-1 DOWNTO 0); 

signal b_xl: std_logic_vector((NB-1)+3 downto 0);

signal partial: pptype;

signal p_0: p_layer_6; -- Top layer
signal p_1: p_layer_5; 
signal p_2: p_layer_4;
signal p_3: p_layer_3;
signal p_4: p_layer_2;
signal p_5: p_layer_1;
signal p_6: p_layer_0;

BEGIN

b_xl(0) <= '0';

b_xl(NB+2 downto NB+1) <= "00";

b_xl(NB downto 1) <= b;


MBEx: for i in 0 to (NB/2 + 1) - 1 generate

		MBE_x0 : MBE
			GENERIC MAP ( NB )
			PORT MAP( a, b_xl(2*i+2 downto 2*i), partial(i));
	
end generate MBEx;


p_0(0)(NB downto 0) <= partial(0);

p_0(0)(NB+3 downto NB+1) <= not(b(1)) & b(1) & b(1);

p_0(1)(0) <= b(1);


tree: for i in 1 to (NB/2 + 1) - 1 - 2 generate

	p_0(i+1)(2*i) <= b(2*i+1);
	
	p_0(i)(NB+2*i downto 2*i) <= partial(i);
	
	p_0(i)(NB+2+2*i downto NB+1+2*i) <= '1' & not(b(2*i+1));

end generate tree;

	
p_0(NB/2-1)(2*NB-2 downto NB-2) <= partial(NB/2-1);

p_0(NB/2-1)(2*NB-1) <= not(b(NB-1));

p_0(NB/2)(NB-2) <= b(NB-1);

p_0(NB/2)(2*NB-1 downto NB) <= partial(NB/2)(NB-1 downto 0);

p_6(1)(1) <= '0';


KS: ks_adder 
	GENERIC MAP(64)
	PORT MAP( a => p_6(0)(2*NB-1 downto 0), b => p_6(1)(2*NB-1 downto 0), sum => prod);

p_1(0)(0) <= p_0(0)(0); 
p_1(0)(1) <= p_0(0)(1); 
p_1(0)(2) <= p_0(0)(2); 
p_1(0)(3) <= p_0(0)(3); 
p_1(0)(4) <= p_0(0)(4); 
p_1(0)(5) <= p_0(0)(5); 
p_1(0)(6) <= p_0(0)(6); 
p_1(0)(7) <= p_0(0)(7); 
p_1(0)(8) <= p_0(0)(8); 
p_1(0)(9) <= p_0(0)(9); 
p_1(0)(10) <= p_0(0)(10); 
p_1(0)(11) <= p_0(0)(11); 
p_1(0)(12) <= p_0(0)(12); 
p_1(0)(13) <= p_0(0)(13); 
p_1(0)(14) <= p_0(0)(14); 
p_1(0)(15) <= p_0(0)(15); 
p_1(0)(16) <= p_0(0)(16); 
p_1(0)(17) <= p_0(0)(17); 
p_1(0)(18) <= p_0(0)(18); 
p_1(0)(19) <= p_0(0)(19); 
p_1(0)(20) <= p_0(0)(20); 
p_1(0)(21) <= p_0(0)(21); 
p_1(0)(22) <= p_0(0)(22); 
p_1(0)(23) <= p_0(0)(23); 
ha_0_24_0: Half_Adder port map( a => p_0(0)(24), b => p_0(1)(24), cout => p_1(12)(25), s => p_1(0)(24)); 
ha_0_25_0: Half_Adder port map( a => p_0(0)(25), b => p_0(1)(25), cout => p_1(12)(26), s => p_1(0)(25)); 
ha_0_26_0: Half_Adder port map( a => p_0(0)(26), b => p_0(1)(26), cout => p_1(12)(27), s => p_1(0)(26)); 
ha_0_27_0: Half_Adder port map( a => p_0(0)(27), b => p_0(1)(27), cout => p_1(12)(28), s => p_1(0)(27)); 
ha_0_28_0: Half_Adder port map( a => p_0(0)(28), b => p_0(1)(28), cout => p_1(12)(29), s => p_1(0)(28)); 
ha_0_29_0: Half_Adder port map( a => p_0(0)(29), b => p_0(1)(29), cout => p_1(12)(30), s => p_1(0)(29)); 
ha_0_30_0: Half_Adder port map( a => p_0(0)(30), b => p_0(1)(30), cout => p_1(12)(31), s => p_1(0)(30)); 
ha_0_31_0: Half_Adder port map( a => p_0(0)(31), b => p_0(1)(31), cout => p_1(12)(32), s => p_1(0)(31)); 
fa_0_32_0: Full_Adder port map( a => p_0(0)(32), b => p_0(1)(32), cin => p_0(2)(32), cout => p_1(12)(33), s => p_1(0)(32)); 
fa_0_33_0: Full_Adder port map( a => p_0(0)(33), b => p_0(1)(33), cin => p_0(2)(33), cout => p_1(12)(34), s => p_1(0)(33)); 
fa_0_34_0: Full_Adder port map( a => p_0(0)(34), b => p_0(1)(34), cin => p_0(2)(34), cout => p_1(12)(35), s => p_1(0)(34)); 
fa_0_35_0: Full_Adder port map( a => p_0(0)(35), b => p_0(1)(35), cin => p_0(2)(35), cout => p_1(12)(36), s => p_1(0)(35)); 
p_1(1)(0) <= p_0(1)(0); 
p_1(1)(2) <= p_0(1)(2); 
p_1(1)(3) <= p_0(1)(3); 
p_1(1)(4) <= p_0(1)(4); 
p_1(1)(5) <= p_0(1)(5); 
p_1(1)(6) <= p_0(1)(6); 
p_1(1)(7) <= p_0(1)(7); 
p_1(1)(8) <= p_0(1)(8); 
p_1(1)(9) <= p_0(1)(9); 
p_1(1)(10) <= p_0(1)(10); 
p_1(1)(11) <= p_0(1)(11); 
p_1(1)(12) <= p_0(1)(12); 
p_1(1)(13) <= p_0(1)(13); 
p_1(1)(14) <= p_0(1)(14); 
p_1(1)(15) <= p_0(1)(15); 
p_1(1)(16) <= p_0(1)(16); 
p_1(1)(17) <= p_0(1)(17); 
p_1(1)(18) <= p_0(1)(18); 
p_1(1)(19) <= p_0(1)(19); 
p_1(1)(20) <= p_0(1)(20); 
p_1(1)(21) <= p_0(1)(21); 
p_1(1)(22) <= p_0(1)(22); 
p_1(1)(23) <= p_0(1)(23); 
ha_0_36_0: Half_Adder port map( a => p_0(1)(36), b => p_0(2)(36), cout => p_1(12)(37), s => p_1(0)(36)); 
p_1(2)(2) <= p_0(2)(2); 
p_1(2)(4) <= p_0(2)(4); 
p_1(2)(5) <= p_0(2)(5); 
p_1(2)(6) <= p_0(2)(6); 
p_1(2)(7) <= p_0(2)(7); 
p_1(2)(8) <= p_0(2)(8); 
p_1(2)(9) <= p_0(2)(9); 
p_1(2)(10) <= p_0(2)(10); 
p_1(2)(11) <= p_0(2)(11); 
p_1(2)(12) <= p_0(2)(12); 
p_1(2)(13) <= p_0(2)(13); 
p_1(2)(14) <= p_0(2)(14); 
p_1(2)(15) <= p_0(2)(15); 
p_1(2)(16) <= p_0(2)(16); 
p_1(2)(17) <= p_0(2)(17); 
p_1(2)(18) <= p_0(2)(18); 
p_1(2)(19) <= p_0(2)(19); 
p_1(2)(20) <= p_0(2)(20); 
p_1(2)(21) <= p_0(2)(21); 
p_1(2)(22) <= p_0(2)(22); 
p_1(2)(23) <= p_0(2)(23); 
p_1(1)(24) <= p_0(2)(24); 
p_1(1)(25) <= p_0(2)(25); 
fa_0_26_0: Full_Adder port map( a => p_0(2)(26), b => p_0(3)(26), cin => p_0(4)(26), cout => p_1(11)(27), s => p_1(1)(26)); 
fa_0_27_0: Full_Adder port map( a => p_0(2)(27), b => p_0(3)(27), cin => p_0(4)(27), cout => p_1(11)(28), s => p_1(1)(27)); 
fa_0_28_0: Full_Adder port map( a => p_0(2)(28), b => p_0(3)(28), cin => p_0(4)(28), cout => p_1(11)(29), s => p_1(1)(28)); 
fa_0_29_0: Full_Adder port map( a => p_0(2)(29), b => p_0(3)(29), cin => p_0(4)(29), cout => p_1(11)(30), s => p_1(1)(29)); 
fa_0_30_0: Full_Adder port map( a => p_0(2)(30), b => p_0(3)(30), cin => p_0(4)(30), cout => p_1(11)(31), s => p_1(1)(30)); 
fa_0_31_0: Full_Adder port map( a => p_0(2)(31), b => p_0(3)(31), cin => p_0(4)(31), cout => p_1(11)(32), s => p_1(1)(31)); 
fa_0_37_0: Full_Adder port map( a => p_0(2)(37), b => p_0(3)(37), cin => p_0(4)(37), cout => p_1(12)(38), s => p_1(0)(37)); 
ha_0_38_0: Half_Adder port map( a => p_0(2)(38), b => p_0(3)(38), cout => p_1(12)(39), s => p_1(0)(38)); 
p_1(3)(4) <= p_0(3)(4); 
p_1(3)(6) <= p_0(3)(6); 
p_1(3)(7) <= p_0(3)(7); 
p_1(3)(8) <= p_0(3)(8); 
p_1(3)(9) <= p_0(3)(9); 
p_1(3)(10) <= p_0(3)(10); 
p_1(3)(11) <= p_0(3)(11); 
p_1(3)(12) <= p_0(3)(12); 
p_1(3)(13) <= p_0(3)(13); 
p_1(3)(14) <= p_0(3)(14); 
p_1(3)(15) <= p_0(3)(15); 
p_1(3)(16) <= p_0(3)(16); 
p_1(3)(17) <= p_0(3)(17); 
p_1(3)(18) <= p_0(3)(18); 
p_1(3)(19) <= p_0(3)(19); 
p_1(3)(20) <= p_0(3)(20); 
p_1(3)(21) <= p_0(3)(21); 
p_1(3)(22) <= p_0(3)(22); 
p_1(3)(23) <= p_0(3)(23); 
p_1(2)(24) <= p_0(3)(24); 
p_1(2)(25) <= p_0(3)(25); 
fa_0_32_1: Full_Adder port map( a => p_0(3)(32), b => p_0(4)(32), cin => p_0(5)(32), cout => p_1(11)(33), s => p_1(1)(32)); 
fa_0_33_1: Full_Adder port map( a => p_0(3)(33), b => p_0(4)(33), cin => p_0(5)(33), cout => p_1(11)(34), s => p_1(1)(33)); 
fa_0_34_1: Full_Adder port map( a => p_0(3)(34), b => p_0(4)(34), cin => p_0(5)(34), cout => p_1(11)(35), s => p_1(1)(34)); 
fa_0_35_1: Full_Adder port map( a => p_0(3)(35), b => p_0(4)(35), cin => p_0(5)(35), cout => p_1(11)(36), s => p_1(1)(35)); 
fa_0_36_0: Full_Adder port map( a => p_0(3)(36), b => p_0(4)(36), cin => p_0(5)(36), cout => p_1(11)(37), s => p_1(1)(36)); 
fa_0_39_0: Full_Adder port map( a => p_0(3)(39), b => p_0(4)(39), cin => p_0(5)(39), cout => p_1(12)(40), s => p_1(0)(39)); 
ha_0_40_0: Half_Adder port map( a => p_0(3)(40), b => p_0(4)(40), cout => p_1(12)(41), s => p_1(0)(40)); 
p_1(4)(6) <= p_0(4)(6); 
p_1(4)(8) <= p_0(4)(8); 
p_1(4)(9) <= p_0(4)(9); 
p_1(4)(10) <= p_0(4)(10); 
p_1(4)(11) <= p_0(4)(11); 
p_1(4)(12) <= p_0(4)(12); 
p_1(4)(13) <= p_0(4)(13); 
p_1(4)(14) <= p_0(4)(14); 
p_1(4)(15) <= p_0(4)(15); 
p_1(4)(16) <= p_0(4)(16); 
p_1(4)(17) <= p_0(4)(17); 
p_1(4)(18) <= p_0(4)(18); 
p_1(4)(19) <= p_0(4)(19); 
p_1(4)(20) <= p_0(4)(20); 
p_1(4)(21) <= p_0(4)(21); 
p_1(4)(22) <= p_0(4)(22); 
p_1(4)(23) <= p_0(4)(23); 
p_1(3)(24) <= p_0(4)(24); 
p_1(3)(25) <= p_0(4)(25); 
fa_0_38_0: Full_Adder port map( a => p_0(4)(38), b => p_0(5)(38), cin => p_0(6)(38), cout => p_1(11)(39), s => p_1(1)(38)); 
fa_0_41_0: Full_Adder port map( a => p_0(4)(41), b => p_0(5)(41), cin => p_0(6)(41), cout => p_1(12)(42), s => p_1(0)(41)); 
ha_0_42_0: Half_Adder port map( a => p_0(4)(42), b => p_0(5)(42), cout => p_1(12)(43), s => p_1(0)(42)); 
p_1(5)(8) <= p_0(5)(8); 
p_1(5)(10) <= p_0(5)(10); 
p_1(5)(11) <= p_0(5)(11); 
p_1(5)(12) <= p_0(5)(12); 
p_1(5)(13) <= p_0(5)(13); 
p_1(5)(14) <= p_0(5)(14); 
p_1(5)(15) <= p_0(5)(15); 
p_1(5)(16) <= p_0(5)(16); 
p_1(5)(17) <= p_0(5)(17); 
p_1(5)(18) <= p_0(5)(18); 
p_1(5)(19) <= p_0(5)(19); 
p_1(5)(20) <= p_0(5)(20); 
p_1(5)(21) <= p_0(5)(21); 
p_1(5)(22) <= p_0(5)(22); 
p_1(5)(23) <= p_0(5)(23); 
p_1(4)(24) <= p_0(5)(24); 
p_1(4)(25) <= p_0(5)(25); 
p_1(2)(26) <= p_0(5)(26); 
p_1(2)(27) <= p_0(5)(27); 
fa_0_28_1: Full_Adder port map( a => p_0(5)(28), b => p_0(6)(28), cin => p_0(7)(28), cout => p_1(10)(29), s => p_1(2)(28)); 
fa_0_29_1: Full_Adder port map( a => p_0(5)(29), b => p_0(6)(29), cin => p_0(7)(29), cout => p_1(10)(30), s => p_1(2)(29)); 
fa_0_30_1: Full_Adder port map( a => p_0(5)(30), b => p_0(6)(30), cin => p_0(7)(30), cout => p_1(10)(31), s => p_1(2)(30)); 
fa_0_31_1: Full_Adder port map( a => p_0(5)(31), b => p_0(6)(31), cin => p_0(7)(31), cout => p_1(10)(32), s => p_1(2)(31)); 
fa_0_37_1: Full_Adder port map( a => p_0(5)(37), b => p_0(6)(37), cin => p_0(7)(37), cout => p_1(11)(38), s => p_1(1)(37)); 
fa_0_40_0: Full_Adder port map( a => p_0(5)(40), b => p_0(6)(40), cin => p_0(7)(40), cout => p_1(11)(41), s => p_1(1)(40)); 
p_1(0)(43) <= p_0(5)(43); 
p_1(0)(44) <= p_0(5)(44); 
p_1(6)(10) <= p_0(6)(10); 
p_1(6)(12) <= p_0(6)(12); 
p_1(6)(13) <= p_0(6)(13); 
p_1(6)(14) <= p_0(6)(14); 
p_1(6)(15) <= p_0(6)(15); 
p_1(6)(16) <= p_0(6)(16); 
p_1(6)(17) <= p_0(6)(17); 
p_1(6)(18) <= p_0(6)(18); 
p_1(6)(19) <= p_0(6)(19); 
p_1(6)(20) <= p_0(6)(20); 
p_1(6)(21) <= p_0(6)(21); 
p_1(6)(22) <= p_0(6)(22); 
p_1(6)(23) <= p_0(6)(23); 
p_1(5)(24) <= p_0(6)(24); 
p_1(5)(25) <= p_0(6)(25); 
p_1(3)(26) <= p_0(6)(26); 
p_1(3)(27) <= p_0(6)(27); 
fa_0_32_2: Full_Adder port map( a => p_0(6)(32), b => p_0(7)(32), cin => p_0(8)(32), cout => p_1(10)(33), s => p_1(2)(32)); 
fa_0_33_2: Full_Adder port map( a => p_0(6)(33), b => p_0(7)(33), cin => p_0(8)(33), cout => p_1(10)(34), s => p_1(2)(33)); 
fa_0_34_2: Full_Adder port map( a => p_0(6)(34), b => p_0(7)(34), cin => p_0(8)(34), cout => p_1(10)(35), s => p_1(2)(34)); 
fa_0_35_2: Full_Adder port map( a => p_0(6)(35), b => p_0(7)(35), cin => p_0(8)(35), cout => p_1(10)(36), s => p_1(2)(35)); 
fa_0_36_1: Full_Adder port map( a => p_0(6)(36), b => p_0(7)(36), cin => p_0(8)(36), cout => p_1(10)(37), s => p_1(2)(36)); 
fa_0_39_1: Full_Adder port map( a => p_0(6)(39), b => p_0(7)(39), cin => p_0(8)(39), cout => p_1(11)(40), s => p_1(1)(39)); 
p_1(1)(42) <= p_0(6)(42); 
p_1(1)(43) <= p_0(6)(43); 
p_1(1)(44) <= p_0(6)(44); 
p_1(0)(45) <= p_0(6)(45); 
p_1(0)(46) <= p_0(6)(46); 
p_1(7)(12) <= p_0(7)(12); 
p_1(7)(14) <= p_0(7)(14); 
p_1(7)(15) <= p_0(7)(15); 
p_1(7)(16) <= p_0(7)(16); 
p_1(7)(17) <= p_0(7)(17); 
p_1(7)(18) <= p_0(7)(18); 
p_1(7)(19) <= p_0(7)(19); 
p_1(7)(20) <= p_0(7)(20); 
p_1(7)(21) <= p_0(7)(21); 
p_1(7)(22) <= p_0(7)(22); 
p_1(7)(23) <= p_0(7)(23); 
p_1(6)(24) <= p_0(7)(24); 
p_1(6)(25) <= p_0(7)(25); 
p_1(4)(26) <= p_0(7)(26); 
p_1(4)(27) <= p_0(7)(27); 
fa_0_38_1: Full_Adder port map( a => p_0(7)(38), b => p_0(8)(38), cin => p_0(9)(38), cout => p_1(10)(39), s => p_1(2)(38)); 
p_1(1)(41) <= p_0(7)(41); 
p_1(2)(42) <= p_0(7)(42); 
p_1(2)(43) <= p_0(7)(43); 
p_1(2)(44) <= p_0(7)(44); 
p_1(1)(45) <= p_0(7)(45); 
p_1(1)(46) <= p_0(7)(46); 
p_1(0)(47) <= p_0(7)(47); 
p_1(0)(48) <= p_0(7)(48); 
p_1(8)(14) <= p_0(8)(14); 
p_1(8)(16) <= p_0(8)(16); 
p_1(8)(17) <= p_0(8)(17); 
p_1(8)(18) <= p_0(8)(18); 
p_1(8)(19) <= p_0(8)(19); 
p_1(8)(20) <= p_0(8)(20); 
p_1(8)(21) <= p_0(8)(21); 
p_1(8)(22) <= p_0(8)(22); 
p_1(8)(23) <= p_0(8)(23); 
p_1(7)(24) <= p_0(8)(24); 
p_1(7)(25) <= p_0(8)(25); 
p_1(5)(26) <= p_0(8)(26); 
p_1(5)(27) <= p_0(8)(27); 
p_1(3)(28) <= p_0(8)(28); 
p_1(3)(29) <= p_0(8)(29); 
fa_0_30_2: Full_Adder port map( a => p_0(8)(30), b => p_0(9)(30), cin => p_0(10)(30), cout => p_1(9)(31), s => p_1(3)(30)); 
fa_0_31_2: Full_Adder port map( a => p_0(8)(31), b => p_0(9)(31), cin => p_0(10)(31), cout => p_1(9)(32), s => p_1(3)(31)); 
fa_0_37_2: Full_Adder port map( a => p_0(8)(37), b => p_0(9)(37), cin => p_0(10)(37), cout => p_1(10)(38), s => p_1(2)(37)); 
p_1(2)(40) <= p_0(8)(40); 
p_1(2)(41) <= p_0(8)(41); 
p_1(3)(42) <= p_0(8)(42); 
p_1(3)(43) <= p_0(8)(43); 
p_1(3)(44) <= p_0(8)(44); 
p_1(2)(45) <= p_0(8)(45); 
p_1(2)(46) <= p_0(8)(46); 
p_1(1)(47) <= p_0(8)(47); 
p_1(1)(48) <= p_0(8)(48); 
p_1(0)(49) <= p_0(8)(49); 
p_1(0)(50) <= p_0(8)(50); 
p_1(9)(16) <= p_0(9)(16); 
p_1(9)(18) <= p_0(9)(18); 
p_1(9)(19) <= p_0(9)(19); 
p_1(9)(20) <= p_0(9)(20); 
p_1(9)(21) <= p_0(9)(21); 
p_1(9)(22) <= p_0(9)(22); 
p_1(9)(23) <= p_0(9)(23); 
p_1(8)(24) <= p_0(9)(24); 
p_1(8)(25) <= p_0(9)(25); 
p_1(6)(26) <= p_0(9)(26); 
p_1(6)(27) <= p_0(9)(27); 
p_1(4)(28) <= p_0(9)(28); 
p_1(4)(29) <= p_0(9)(29); 
fa_0_32_3: Full_Adder port map( a => p_0(9)(32), b => p_0(10)(32), cin => p_0(11)(32), cout => p_1(9)(33), s => p_1(3)(32)); 
fa_0_33_3: Full_Adder port map( a => p_0(9)(33), b => p_0(10)(33), cin => p_0(11)(33), cout => p_1(9)(34), s => p_1(3)(33)); 
fa_0_34_3: Full_Adder port map( a => p_0(9)(34), b => p_0(10)(34), cin => p_0(11)(34), cout => p_1(9)(35), s => p_1(3)(34)); 
fa_0_35_3: Full_Adder port map( a => p_0(9)(35), b => p_0(10)(35), cin => p_0(11)(35), cout => p_1(9)(36), s => p_1(3)(35)); 
fa_0_36_2: Full_Adder port map( a => p_0(9)(36), b => p_0(10)(36), cin => p_0(11)(36), cout => p_1(9)(37), s => p_1(3)(36)); 
p_1(2)(39) <= p_0(9)(39); 
p_1(3)(40) <= p_0(9)(40); 
p_1(3)(41) <= p_0(9)(41); 
p_1(4)(42) <= p_0(9)(42); 
p_1(4)(43) <= p_0(9)(43); 
p_1(4)(44) <= p_0(9)(44); 
p_1(3)(45) <= p_0(9)(45); 
p_1(3)(46) <= p_0(9)(46); 
p_1(2)(47) <= p_0(9)(47); 
p_1(2)(48) <= p_0(9)(48); 
p_1(1)(49) <= p_0(9)(49); 
p_1(1)(50) <= p_0(9)(50); 
p_1(0)(51) <= p_0(9)(51); 
p_1(0)(52) <= p_0(9)(52); 
p_1(10)(18) <= p_0(10)(18); 
p_1(10)(20) <= p_0(10)(20); 
p_1(10)(21) <= p_0(10)(21); 
p_1(10)(22) <= p_0(10)(22); 
p_1(10)(23) <= p_0(10)(23); 
p_1(9)(24) <= p_0(10)(24); 
p_1(9)(25) <= p_0(10)(25); 
p_1(7)(26) <= p_0(10)(26); 
p_1(7)(27) <= p_0(10)(27); 
p_1(5)(28) <= p_0(10)(28); 
p_1(5)(29) <= p_0(10)(29); 
p_1(3)(38) <= p_0(10)(38); 
p_1(3)(39) <= p_0(10)(39); 
p_1(4)(40) <= p_0(10)(40); 
p_1(4)(41) <= p_0(10)(41); 
p_1(5)(42) <= p_0(10)(42); 
p_1(5)(43) <= p_0(10)(43); 
p_1(5)(44) <= p_0(10)(44); 
p_1(4)(45) <= p_0(10)(45); 
p_1(4)(46) <= p_0(10)(46); 
p_1(3)(47) <= p_0(10)(47); 
p_1(3)(48) <= p_0(10)(48); 
p_1(2)(49) <= p_0(10)(49); 
p_1(2)(50) <= p_0(10)(50); 
p_1(1)(51) <= p_0(10)(51); 
p_1(1)(52) <= p_0(10)(52); 
p_1(0)(53) <= p_0(10)(53); 
p_1(0)(54) <= p_0(10)(54); 
p_1(11)(20) <= p_0(11)(20); 
p_1(11)(22) <= p_0(11)(22); 
p_1(11)(23) <= p_0(11)(23); 
p_1(10)(24) <= p_0(11)(24); 
p_1(10)(25) <= p_0(11)(25); 
p_1(8)(26) <= p_0(11)(26); 
p_1(8)(27) <= p_0(11)(27); 
p_1(6)(28) <= p_0(11)(28); 
p_1(6)(29) <= p_0(11)(29); 
p_1(4)(30) <= p_0(11)(30); 
p_1(4)(31) <= p_0(11)(31); 
p_1(3)(37) <= p_0(11)(37); 
p_1(4)(38) <= p_0(11)(38); 
p_1(4)(39) <= p_0(11)(39); 
p_1(5)(40) <= p_0(11)(40); 
p_1(5)(41) <= p_0(11)(41); 
p_1(6)(42) <= p_0(11)(42); 
p_1(6)(43) <= p_0(11)(43); 
p_1(6)(44) <= p_0(11)(44); 
p_1(5)(45) <= p_0(11)(45); 
p_1(5)(46) <= p_0(11)(46); 
p_1(4)(47) <= p_0(11)(47); 
p_1(4)(48) <= p_0(11)(48); 
p_1(3)(49) <= p_0(11)(49); 
p_1(3)(50) <= p_0(11)(50); 
p_1(2)(51) <= p_0(11)(51); 
p_1(2)(52) <= p_0(11)(52); 
p_1(1)(53) <= p_0(11)(53); 
p_1(1)(54) <= p_0(11)(54); 
p_1(0)(55) <= p_0(11)(55); 
p_1(0)(56) <= p_0(11)(56); 
p_1(12)(22) <= p_0(12)(22); 
p_1(11)(24) <= p_0(12)(24); 
p_1(11)(25) <= p_0(12)(25); 
p_1(9)(26) <= p_0(12)(26); 
p_1(9)(27) <= p_0(12)(27); 
p_1(7)(28) <= p_0(12)(28); 
p_1(7)(29) <= p_0(12)(29); 
p_1(5)(30) <= p_0(12)(30); 
p_1(5)(31) <= p_0(12)(31); 
p_1(4)(32) <= p_0(12)(32); 
p_1(4)(33) <= p_0(12)(33); 
p_1(4)(34) <= p_0(12)(34); 
p_1(4)(35) <= p_0(12)(35); 
p_1(4)(36) <= p_0(12)(36); 
p_1(4)(37) <= p_0(12)(37); 
p_1(5)(38) <= p_0(12)(38); 
p_1(5)(39) <= p_0(12)(39); 
p_1(6)(40) <= p_0(12)(40); 
p_1(6)(41) <= p_0(12)(41); 
p_1(7)(42) <= p_0(12)(42); 
p_1(7)(43) <= p_0(12)(43); 
p_1(7)(44) <= p_0(12)(44); 
p_1(6)(45) <= p_0(12)(45); 
p_1(6)(46) <= p_0(12)(46); 
p_1(5)(47) <= p_0(12)(47); 
p_1(5)(48) <= p_0(12)(48); 
p_1(4)(49) <= p_0(12)(49); 
p_1(4)(50) <= p_0(12)(50); 
p_1(3)(51) <= p_0(12)(51); 
p_1(3)(52) <= p_0(12)(52); 
p_1(2)(53) <= p_0(12)(53); 
p_1(2)(54) <= p_0(12)(54); 
p_1(1)(55) <= p_0(12)(55); 
p_1(1)(56) <= p_0(12)(56); 
p_1(0)(57) <= p_0(12)(57); 
p_1(0)(58) <= p_0(12)(58); 
p_1(12)(24) <= p_0(13)(24); 
p_1(10)(26) <= p_0(13)(26); 
p_1(10)(27) <= p_0(13)(27); 
p_1(8)(28) <= p_0(13)(28); 
p_1(8)(29) <= p_0(13)(29); 
p_1(6)(30) <= p_0(13)(30); 
p_1(6)(31) <= p_0(13)(31); 
p_1(5)(32) <= p_0(13)(32); 
p_1(5)(33) <= p_0(13)(33); 
p_1(5)(34) <= p_0(13)(34); 
p_1(5)(35) <= p_0(13)(35); 
p_1(5)(36) <= p_0(13)(36); 
p_1(5)(37) <= p_0(13)(37); 
p_1(6)(38) <= p_0(13)(38); 
p_1(6)(39) <= p_0(13)(39); 
p_1(7)(40) <= p_0(13)(40); 
p_1(7)(41) <= p_0(13)(41); 
p_1(8)(42) <= p_0(13)(42); 
p_1(8)(43) <= p_0(13)(43); 
p_1(8)(44) <= p_0(13)(44); 
p_1(7)(45) <= p_0(13)(45); 
p_1(7)(46) <= p_0(13)(46); 
p_1(6)(47) <= p_0(13)(47); 
p_1(6)(48) <= p_0(13)(48); 
p_1(5)(49) <= p_0(13)(49); 
p_1(5)(50) <= p_0(13)(50); 
p_1(4)(51) <= p_0(13)(51); 
p_1(4)(52) <= p_0(13)(52); 
p_1(3)(53) <= p_0(13)(53); 
p_1(3)(54) <= p_0(13)(54); 
p_1(2)(55) <= p_0(13)(55); 
p_1(2)(56) <= p_0(13)(56); 
p_1(1)(57) <= p_0(13)(57); 
p_1(1)(58) <= p_0(13)(58); 
p_1(0)(59) <= p_0(13)(59); 
p_1(0)(60) <= p_0(13)(60); 
p_1(11)(26) <= p_0(14)(26); 
p_1(9)(28) <= p_0(14)(28); 
p_1(9)(29) <= p_0(14)(29); 
p_1(7)(30) <= p_0(14)(30); 
p_1(7)(31) <= p_0(14)(31); 
p_1(6)(32) <= p_0(14)(32); 
p_1(6)(33) <= p_0(14)(33); 
p_1(6)(34) <= p_0(14)(34); 
p_1(6)(35) <= p_0(14)(35); 
p_1(6)(36) <= p_0(14)(36); 
p_1(6)(37) <= p_0(14)(37); 
p_1(7)(38) <= p_0(14)(38); 
p_1(7)(39) <= p_0(14)(39); 
p_1(8)(40) <= p_0(14)(40); 
p_1(8)(41) <= p_0(14)(41); 
p_1(9)(42) <= p_0(14)(42); 
p_1(9)(43) <= p_0(14)(43); 
p_1(9)(44) <= p_0(14)(44); 
p_1(8)(45) <= p_0(14)(45); 
p_1(8)(46) <= p_0(14)(46); 
p_1(7)(47) <= p_0(14)(47); 
p_1(7)(48) <= p_0(14)(48); 
p_1(6)(49) <= p_0(14)(49); 
p_1(6)(50) <= p_0(14)(50); 
p_1(5)(51) <= p_0(14)(51); 
p_1(5)(52) <= p_0(14)(52); 
p_1(4)(53) <= p_0(14)(53); 
p_1(4)(54) <= p_0(14)(54); 
p_1(3)(55) <= p_0(14)(55); 
p_1(3)(56) <= p_0(14)(56); 
p_1(2)(57) <= p_0(14)(57); 
p_1(2)(58) <= p_0(14)(58); 
p_1(1)(59) <= p_0(14)(59); 
p_1(1)(60) <= p_0(14)(60); 
p_1(0)(61) <= p_0(14)(61); 
p_1(0)(62) <= p_0(14)(62); 
p_1(10)(28) <= p_0(15)(28); 
p_1(8)(30) <= p_0(15)(30); 
p_1(8)(31) <= p_0(15)(31); 
p_1(7)(32) <= p_0(15)(32); 
p_1(7)(33) <= p_0(15)(33); 
p_1(7)(34) <= p_0(15)(34); 
p_1(7)(35) <= p_0(15)(35); 
p_1(7)(36) <= p_0(15)(36); 
p_1(7)(37) <= p_0(15)(37); 
p_1(8)(38) <= p_0(15)(38); 
p_1(8)(39) <= p_0(15)(39); 
p_1(9)(40) <= p_0(15)(40); 
p_1(9)(41) <= p_0(15)(41); 
p_1(10)(42) <= p_0(15)(42); 
p_1(10)(43) <= p_0(15)(43); 
p_1(10)(44) <= p_0(15)(44); 
p_1(9)(45) <= p_0(15)(45); 
p_1(9)(46) <= p_0(15)(46); 
p_1(8)(47) <= p_0(15)(47); 
p_1(8)(48) <= p_0(15)(48); 
p_1(7)(49) <= p_0(15)(49); 
p_1(7)(50) <= p_0(15)(50); 
p_1(6)(51) <= p_0(15)(51); 
p_1(6)(52) <= p_0(15)(52); 
p_1(5)(53) <= p_0(15)(53); 
p_1(5)(54) <= p_0(15)(54); 
p_1(4)(55) <= p_0(15)(55); 
p_1(4)(56) <= p_0(15)(56); 
p_1(3)(57) <= p_0(15)(57); 
p_1(3)(58) <= p_0(15)(58); 
p_1(2)(59) <= p_0(15)(59); 
p_1(2)(60) <= p_0(15)(60); 
p_1(1)(61) <= p_0(15)(61); 
p_1(1)(62) <= p_0(15)(62); 
p_1(0)(63) <= p_0(15)(63); 
p_1(9)(30) <= p_0(16)(30); 
p_1(8)(32) <= p_0(16)(32); 
p_1(8)(33) <= p_0(16)(33); 
p_1(8)(34) <= p_0(16)(34); 
p_1(8)(35) <= p_0(16)(35); 
p_1(8)(36) <= p_0(16)(36); 
p_1(8)(37) <= p_0(16)(37); 
p_1(9)(38) <= p_0(16)(38); 
p_1(9)(39) <= p_0(16)(39); 
p_1(10)(40) <= p_0(16)(40); 
p_1(10)(41) <= p_0(16)(41); 
p_1(11)(42) <= p_0(16)(42); 
p_1(11)(43) <= p_0(16)(43); 
p_1(11)(44) <= p_0(16)(44); 
p_1(10)(45) <= p_0(16)(45); 
p_1(10)(46) <= p_0(16)(46); 
p_1(9)(47) <= p_0(16)(47); 
p_1(9)(48) <= p_0(16)(48); 
p_1(8)(49) <= p_0(16)(49); 
p_1(8)(50) <= p_0(16)(50); 
p_1(7)(51) <= p_0(16)(51); 
p_1(7)(52) <= p_0(16)(52); 
p_1(6)(53) <= p_0(16)(53); 
p_1(6)(54) <= p_0(16)(54); 
p_1(5)(55) <= p_0(16)(55); 
p_1(5)(56) <= p_0(16)(56); 
p_1(4)(57) <= p_0(16)(57); 
p_1(4)(58) <= p_0(16)(58); 
p_1(3)(59) <= p_0(16)(59); 
p_1(3)(60) <= p_0(16)(60); 
p_1(2)(61) <= p_0(16)(61); 
p_1(2)(62) <= p_0(16)(62); 
p_1(1)(63) <= p_0(16)(63); 
p_2(0)(0) <= p_1(0)(0); 
p_2(0)(1) <= p_1(0)(1); 
p_2(0)(2) <= p_1(0)(2); 
p_2(0)(3) <= p_1(0)(3); 
p_2(0)(4) <= p_1(0)(4); 
p_2(0)(5) <= p_1(0)(5); 
p_2(0)(6) <= p_1(0)(6); 
p_2(0)(7) <= p_1(0)(7); 
p_2(0)(8) <= p_1(0)(8); 
p_2(0)(9) <= p_1(0)(9); 
p_2(0)(10) <= p_1(0)(10); 
p_2(0)(11) <= p_1(0)(11); 
p_2(0)(12) <= p_1(0)(12); 
p_2(0)(13) <= p_1(0)(13); 
p_2(0)(14) <= p_1(0)(14); 
p_2(0)(15) <= p_1(0)(15); 
ha_1_16_0: Half_Adder port map( a => p_1(0)(16), b => p_1(1)(16), cout => p_2(8)(17), s => p_2(0)(16)); 
ha_1_17_0: Half_Adder port map( a => p_1(0)(17), b => p_1(1)(17), cout => p_2(8)(18), s => p_2(0)(17)); 
ha_1_18_0: Half_Adder port map( a => p_1(0)(18), b => p_1(1)(18), cout => p_2(8)(19), s => p_2(0)(18)); 
ha_1_19_0: Half_Adder port map( a => p_1(0)(19), b => p_1(1)(19), cout => p_2(8)(20), s => p_2(0)(19)); 
ha_1_20_0: Half_Adder port map( a => p_1(0)(20), b => p_1(1)(20), cout => p_2(8)(21), s => p_2(0)(20)); 
ha_1_21_0: Half_Adder port map( a => p_1(0)(21), b => p_1(1)(21), cout => p_2(8)(22), s => p_2(0)(21)); 
ha_1_22_0: Half_Adder port map( a => p_1(0)(22), b => p_1(1)(22), cout => p_2(8)(23), s => p_2(0)(22)); 
ha_1_23_0: Half_Adder port map( a => p_1(0)(23), b => p_1(1)(23), cout => p_2(8)(24), s => p_2(0)(23)); 
fa_1_24_0: Full_Adder port map( a => p_1(0)(24), b => p_1(1)(24), cin => p_1(2)(24), cout => p_2(8)(25), s => p_2(0)(24)); 
fa_1_25_0: Full_Adder port map( a => p_1(0)(25), b => p_1(1)(25), cin => p_1(2)(25), cout => p_2(8)(26), s => p_2(0)(25)); 
fa_1_26_0: Full_Adder port map( a => p_1(0)(26), b => p_1(1)(26), cin => p_1(2)(26), cout => p_2(8)(27), s => p_2(0)(26)); 
fa_1_27_0: Full_Adder port map( a => p_1(0)(27), b => p_1(1)(27), cin => p_1(2)(27), cout => p_2(8)(28), s => p_2(0)(27)); 
fa_1_28_0: Full_Adder port map( a => p_1(0)(28), b => p_1(1)(28), cin => p_1(2)(28), cout => p_2(8)(29), s => p_2(0)(28)); 
fa_1_29_0: Full_Adder port map( a => p_1(0)(29), b => p_1(1)(29), cin => p_1(2)(29), cout => p_2(8)(30), s => p_2(0)(29)); 
fa_1_30_0: Full_Adder port map( a => p_1(0)(30), b => p_1(1)(30), cin => p_1(2)(30), cout => p_2(8)(31), s => p_2(0)(30)); 
fa_1_31_0: Full_Adder port map( a => p_1(0)(31), b => p_1(1)(31), cin => p_1(2)(31), cout => p_2(8)(32), s => p_2(0)(31)); 
fa_1_32_0: Full_Adder port map( a => p_1(0)(32), b => p_1(1)(32), cin => p_1(2)(32), cout => p_2(8)(33), s => p_2(0)(32)); 
fa_1_33_0: Full_Adder port map( a => p_1(0)(33), b => p_1(1)(33), cin => p_1(2)(33), cout => p_2(8)(34), s => p_2(0)(33)); 
fa_1_34_0: Full_Adder port map( a => p_1(0)(34), b => p_1(1)(34), cin => p_1(2)(34), cout => p_2(8)(35), s => p_2(0)(34)); 
fa_1_35_0: Full_Adder port map( a => p_1(0)(35), b => p_1(1)(35), cin => p_1(2)(35), cout => p_2(8)(36), s => p_2(0)(35)); 
fa_1_36_0: Full_Adder port map( a => p_1(0)(36), b => p_1(1)(36), cin => p_1(2)(36), cout => p_2(8)(37), s => p_2(0)(36)); 
fa_1_37_0: Full_Adder port map( a => p_1(0)(37), b => p_1(1)(37), cin => p_1(2)(37), cout => p_2(8)(38), s => p_2(0)(37)); 
fa_1_38_0: Full_Adder port map( a => p_1(0)(38), b => p_1(1)(38), cin => p_1(2)(38), cout => p_2(8)(39), s => p_2(0)(38)); 
fa_1_39_0: Full_Adder port map( a => p_1(0)(39), b => p_1(1)(39), cin => p_1(2)(39), cout => p_2(8)(40), s => p_2(0)(39)); 
fa_1_40_0: Full_Adder port map( a => p_1(0)(40), b => p_1(1)(40), cin => p_1(2)(40), cout => p_2(8)(41), s => p_2(0)(40)); 
fa_1_41_0: Full_Adder port map( a => p_1(0)(41), b => p_1(1)(41), cin => p_1(2)(41), cout => p_2(8)(42), s => p_2(0)(41)); 
fa_1_42_0: Full_Adder port map( a => p_1(0)(42), b => p_1(1)(42), cin => p_1(2)(42), cout => p_2(8)(43), s => p_2(0)(42)); 
fa_1_43_0: Full_Adder port map( a => p_1(0)(43), b => p_1(1)(43), cin => p_1(2)(43), cout => p_2(8)(44), s => p_2(0)(43)); 
ha_1_44_0: Half_Adder port map( a => p_1(0)(44), b => p_1(1)(44), cout => p_2(8)(45), s => p_2(0)(44)); 
fa_1_45_0: Full_Adder port map( a => p_1(0)(45), b => p_1(1)(45), cin => p_1(2)(45), cout => p_2(8)(46), s => p_2(0)(45)); 
ha_1_46_0: Half_Adder port map( a => p_1(0)(46), b => p_1(1)(46), cout => p_2(8)(47), s => p_2(0)(46)); 
fa_1_47_0: Full_Adder port map( a => p_1(0)(47), b => p_1(1)(47), cin => p_1(2)(47), cout => p_2(8)(48), s => p_2(0)(47)); 
ha_1_48_0: Half_Adder port map( a => p_1(0)(48), b => p_1(1)(48), cout => p_2(8)(49), s => p_2(0)(48)); 
fa_1_49_0: Full_Adder port map( a => p_1(0)(49), b => p_1(1)(49), cin => p_1(2)(49), cout => p_2(8)(50), s => p_2(0)(49)); 
ha_1_50_0: Half_Adder port map( a => p_1(0)(50), b => p_1(1)(50), cout => p_2(8)(51), s => p_2(0)(50)); 
p_2(0)(51) <= p_1(0)(51); 
p_2(0)(52) <= p_1(0)(52); 
p_2(0)(53) <= p_1(0)(53); 
p_2(0)(54) <= p_1(0)(54); 
p_2(0)(55) <= p_1(0)(55); 
p_2(0)(56) <= p_1(0)(56); 
p_2(0)(57) <= p_1(0)(57); 
p_2(0)(58) <= p_1(0)(58); 
p_2(0)(59) <= p_1(0)(59); 
p_2(0)(60) <= p_1(0)(60); 
p_2(0)(61) <= p_1(0)(61); 
p_2(0)(62) <= p_1(0)(62); 
p_2(0)(63) <= p_1(0)(63); 
p_2(1)(0) <= p_1(1)(0); 
p_2(1)(2) <= p_1(1)(2); 
p_2(1)(3) <= p_1(1)(3); 
p_2(1)(4) <= p_1(1)(4); 
p_2(1)(5) <= p_1(1)(5); 
p_2(1)(6) <= p_1(1)(6); 
p_2(1)(7) <= p_1(1)(7); 
p_2(1)(8) <= p_1(1)(8); 
p_2(1)(9) <= p_1(1)(9); 
p_2(1)(10) <= p_1(1)(10); 
p_2(1)(11) <= p_1(1)(11); 
p_2(1)(12) <= p_1(1)(12); 
p_2(1)(13) <= p_1(1)(13); 
p_2(1)(14) <= p_1(1)(14); 
p_2(1)(15) <= p_1(1)(15); 
p_2(1)(51) <= p_1(1)(51); 
p_2(1)(52) <= p_1(1)(52); 
p_2(1)(53) <= p_1(1)(53); 
p_2(1)(54) <= p_1(1)(54); 
p_2(1)(55) <= p_1(1)(55); 
p_2(1)(56) <= p_1(1)(56); 
p_2(1)(57) <= p_1(1)(57); 
p_2(1)(58) <= p_1(1)(58); 
p_2(1)(59) <= p_1(1)(59); 
p_2(1)(60) <= p_1(1)(60); 
p_2(1)(61) <= p_1(1)(61); 
p_2(1)(62) <= p_1(1)(62); 
p_2(1)(63) <= p_1(1)(63); 
p_2(2)(2) <= p_1(2)(2); 
p_2(2)(4) <= p_1(2)(4); 
p_2(2)(5) <= p_1(2)(5); 
p_2(2)(6) <= p_1(2)(6); 
p_2(2)(7) <= p_1(2)(7); 
p_2(2)(8) <= p_1(2)(8); 
p_2(2)(9) <= p_1(2)(9); 
p_2(2)(10) <= p_1(2)(10); 
p_2(2)(11) <= p_1(2)(11); 
p_2(2)(12) <= p_1(2)(12); 
p_2(2)(13) <= p_1(2)(13); 
p_2(2)(14) <= p_1(2)(14); 
p_2(2)(15) <= p_1(2)(15); 
p_2(1)(16) <= p_1(2)(16); 
p_2(1)(17) <= p_1(2)(17); 
fa_1_18_0: Full_Adder port map( a => p_1(2)(18), b => p_1(3)(18), cin => p_1(4)(18), cout => p_2(7)(19), s => p_2(1)(18)); 
fa_1_19_0: Full_Adder port map( a => p_1(2)(19), b => p_1(3)(19), cin => p_1(4)(19), cout => p_2(7)(20), s => p_2(1)(19)); 
fa_1_20_0: Full_Adder port map( a => p_1(2)(20), b => p_1(3)(20), cin => p_1(4)(20), cout => p_2(7)(21), s => p_2(1)(20)); 
fa_1_21_0: Full_Adder port map( a => p_1(2)(21), b => p_1(3)(21), cin => p_1(4)(21), cout => p_2(7)(22), s => p_2(1)(21)); 
fa_1_22_0: Full_Adder port map( a => p_1(2)(22), b => p_1(3)(22), cin => p_1(4)(22), cout => p_2(7)(23), s => p_2(1)(22)); 
fa_1_23_0: Full_Adder port map( a => p_1(2)(23), b => p_1(3)(23), cin => p_1(4)(23), cout => p_2(7)(24), s => p_2(1)(23)); 
fa_1_44_0: Full_Adder port map( a => p_1(2)(44), b => p_1(3)(44), cin => p_1(4)(44), cout => p_2(7)(45), s => p_2(1)(44)); 
fa_1_46_0: Full_Adder port map( a => p_1(2)(46), b => p_1(3)(46), cin => p_1(4)(46), cout => p_2(7)(47), s => p_2(1)(46)); 
fa_1_48_0: Full_Adder port map( a => p_1(2)(48), b => p_1(3)(48), cin => p_1(4)(48), cout => p_2(7)(49), s => p_2(1)(48)); 
p_2(1)(50) <= p_1(2)(50); 
p_2(2)(51) <= p_1(2)(51); 
p_2(2)(52) <= p_1(2)(52); 
p_2(2)(53) <= p_1(2)(53); 
p_2(2)(54) <= p_1(2)(54); 
p_2(2)(55) <= p_1(2)(55); 
p_2(2)(56) <= p_1(2)(56); 
p_2(2)(57) <= p_1(2)(57); 
p_2(2)(58) <= p_1(2)(58); 
p_2(2)(59) <= p_1(2)(59); 
p_2(2)(60) <= p_1(2)(60); 
p_2(2)(61) <= p_1(2)(61); 
p_2(2)(62) <= p_1(2)(62); 
p_2(3)(4) <= p_1(3)(4); 
p_2(3)(6) <= p_1(3)(6); 
p_2(3)(7) <= p_1(3)(7); 
p_2(3)(8) <= p_1(3)(8); 
p_2(3)(9) <= p_1(3)(9); 
p_2(3)(10) <= p_1(3)(10); 
p_2(3)(11) <= p_1(3)(11); 
p_2(3)(12) <= p_1(3)(12); 
p_2(3)(13) <= p_1(3)(13); 
p_2(3)(14) <= p_1(3)(14); 
p_2(3)(15) <= p_1(3)(15); 
p_2(2)(16) <= p_1(3)(16); 
p_2(2)(17) <= p_1(3)(17); 
fa_1_24_1: Full_Adder port map( a => p_1(3)(24), b => p_1(4)(24), cin => p_1(5)(24), cout => p_2(7)(25), s => p_2(1)(24)); 
fa_1_25_1: Full_Adder port map( a => p_1(3)(25), b => p_1(4)(25), cin => p_1(5)(25), cout => p_2(7)(26), s => p_2(1)(25)); 
fa_1_26_1: Full_Adder port map( a => p_1(3)(26), b => p_1(4)(26), cin => p_1(5)(26), cout => p_2(7)(27), s => p_2(1)(26)); 
fa_1_27_1: Full_Adder port map( a => p_1(3)(27), b => p_1(4)(27), cin => p_1(5)(27), cout => p_2(7)(28), s => p_2(1)(27)); 
fa_1_28_1: Full_Adder port map( a => p_1(3)(28), b => p_1(4)(28), cin => p_1(5)(28), cout => p_2(7)(29), s => p_2(1)(28)); 
fa_1_29_1: Full_Adder port map( a => p_1(3)(29), b => p_1(4)(29), cin => p_1(5)(29), cout => p_2(7)(30), s => p_2(1)(29)); 
fa_1_30_1: Full_Adder port map( a => p_1(3)(30), b => p_1(4)(30), cin => p_1(5)(30), cout => p_2(7)(31), s => p_2(1)(30)); 
fa_1_31_1: Full_Adder port map( a => p_1(3)(31), b => p_1(4)(31), cin => p_1(5)(31), cout => p_2(7)(32), s => p_2(1)(31)); 
fa_1_32_1: Full_Adder port map( a => p_1(3)(32), b => p_1(4)(32), cin => p_1(5)(32), cout => p_2(7)(33), s => p_2(1)(32)); 
fa_1_33_1: Full_Adder port map( a => p_1(3)(33), b => p_1(4)(33), cin => p_1(5)(33), cout => p_2(7)(34), s => p_2(1)(33)); 
fa_1_34_1: Full_Adder port map( a => p_1(3)(34), b => p_1(4)(34), cin => p_1(5)(34), cout => p_2(7)(35), s => p_2(1)(34)); 
fa_1_35_1: Full_Adder port map( a => p_1(3)(35), b => p_1(4)(35), cin => p_1(5)(35), cout => p_2(7)(36), s => p_2(1)(35)); 
fa_1_36_1: Full_Adder port map( a => p_1(3)(36), b => p_1(4)(36), cin => p_1(5)(36), cout => p_2(7)(37), s => p_2(1)(36)); 
fa_1_37_1: Full_Adder port map( a => p_1(3)(37), b => p_1(4)(37), cin => p_1(5)(37), cout => p_2(7)(38), s => p_2(1)(37)); 
fa_1_38_1: Full_Adder port map( a => p_1(3)(38), b => p_1(4)(38), cin => p_1(5)(38), cout => p_2(7)(39), s => p_2(1)(38)); 
fa_1_39_1: Full_Adder port map( a => p_1(3)(39), b => p_1(4)(39), cin => p_1(5)(39), cout => p_2(7)(40), s => p_2(1)(39)); 
fa_1_40_1: Full_Adder port map( a => p_1(3)(40), b => p_1(4)(40), cin => p_1(5)(40), cout => p_2(7)(41), s => p_2(1)(40)); 
fa_1_41_1: Full_Adder port map( a => p_1(3)(41), b => p_1(4)(41), cin => p_1(5)(41), cout => p_2(7)(42), s => p_2(1)(41)); 
fa_1_42_1: Full_Adder port map( a => p_1(3)(42), b => p_1(4)(42), cin => p_1(5)(42), cout => p_2(7)(43), s => p_2(1)(42)); 
fa_1_43_1: Full_Adder port map( a => p_1(3)(43), b => p_1(4)(43), cin => p_1(5)(43), cout => p_2(7)(44), s => p_2(1)(43)); 
fa_1_45_1: Full_Adder port map( a => p_1(3)(45), b => p_1(4)(45), cin => p_1(5)(45), cout => p_2(7)(46), s => p_2(1)(45)); 
fa_1_47_1: Full_Adder port map( a => p_1(3)(47), b => p_1(4)(47), cin => p_1(5)(47), cout => p_2(7)(48), s => p_2(1)(47)); 
p_2(1)(49) <= p_1(3)(49); 
p_2(2)(50) <= p_1(3)(50); 
p_2(3)(51) <= p_1(3)(51); 
p_2(3)(52) <= p_1(3)(52); 
p_2(3)(53) <= p_1(3)(53); 
p_2(3)(54) <= p_1(3)(54); 
p_2(3)(55) <= p_1(3)(55); 
p_2(3)(56) <= p_1(3)(56); 
p_2(3)(57) <= p_1(3)(57); 
p_2(3)(58) <= p_1(3)(58); 
p_2(3)(59) <= p_1(3)(59); 
p_2(3)(60) <= p_1(3)(60); 
p_2(4)(6) <= p_1(4)(6); 
p_2(4)(8) <= p_1(4)(8); 
p_2(4)(9) <= p_1(4)(9); 
p_2(4)(10) <= p_1(4)(10); 
p_2(4)(11) <= p_1(4)(11); 
p_2(4)(12) <= p_1(4)(12); 
p_2(4)(13) <= p_1(4)(13); 
p_2(4)(14) <= p_1(4)(14); 
p_2(4)(15) <= p_1(4)(15); 
p_2(3)(16) <= p_1(4)(16); 
p_2(3)(17) <= p_1(4)(17); 
p_2(2)(49) <= p_1(4)(49); 
p_2(3)(50) <= p_1(4)(50); 
p_2(4)(51) <= p_1(4)(51); 
p_2(4)(52) <= p_1(4)(52); 
p_2(4)(53) <= p_1(4)(53); 
p_2(4)(54) <= p_1(4)(54); 
p_2(4)(55) <= p_1(4)(55); 
p_2(4)(56) <= p_1(4)(56); 
p_2(4)(57) <= p_1(4)(57); 
p_2(4)(58) <= p_1(4)(58); 
p_2(5)(8) <= p_1(5)(8); 
p_2(5)(10) <= p_1(5)(10); 
p_2(5)(11) <= p_1(5)(11); 
p_2(5)(12) <= p_1(5)(12); 
p_2(5)(13) <= p_1(5)(13); 
p_2(5)(14) <= p_1(5)(14); 
p_2(5)(15) <= p_1(5)(15); 
p_2(4)(16) <= p_1(5)(16); 
p_2(4)(17) <= p_1(5)(17); 
p_2(2)(18) <= p_1(5)(18); 
p_2(2)(19) <= p_1(5)(19); 
fa_1_20_1: Full_Adder port map( a => p_1(5)(20), b => p_1(6)(20), cin => p_1(7)(20), cout => p_2(6)(21), s => p_2(2)(20)); 
fa_1_21_1: Full_Adder port map( a => p_1(5)(21), b => p_1(6)(21), cin => p_1(7)(21), cout => p_2(6)(22), s => p_2(2)(21)); 
fa_1_22_1: Full_Adder port map( a => p_1(5)(22), b => p_1(6)(22), cin => p_1(7)(22), cout => p_2(6)(23), s => p_2(2)(22)); 
fa_1_23_1: Full_Adder port map( a => p_1(5)(23), b => p_1(6)(23), cin => p_1(7)(23), cout => p_2(6)(24), s => p_2(2)(23)); 
fa_1_44_1: Full_Adder port map( a => p_1(5)(44), b => p_1(6)(44), cin => p_1(7)(44), cout => p_2(6)(45), s => p_2(2)(44)); 
fa_1_46_1: Full_Adder port map( a => p_1(5)(46), b => p_1(6)(46), cin => p_1(7)(46), cout => p_2(6)(47), s => p_2(2)(46)); 
p_2(2)(48) <= p_1(5)(48); 
p_2(3)(49) <= p_1(5)(49); 
p_2(4)(50) <= p_1(5)(50); 
p_2(5)(51) <= p_1(5)(51); 
p_2(5)(52) <= p_1(5)(52); 
p_2(5)(53) <= p_1(5)(53); 
p_2(5)(54) <= p_1(5)(54); 
p_2(5)(55) <= p_1(5)(55); 
p_2(5)(56) <= p_1(5)(56); 
p_2(6)(10) <= p_1(6)(10); 
p_2(6)(12) <= p_1(6)(12); 
p_2(6)(13) <= p_1(6)(13); 
p_2(6)(14) <= p_1(6)(14); 
p_2(6)(15) <= p_1(6)(15); 
p_2(5)(16) <= p_1(6)(16); 
p_2(5)(17) <= p_1(6)(17); 
p_2(3)(18) <= p_1(6)(18); 
p_2(3)(19) <= p_1(6)(19); 
fa_1_24_2: Full_Adder port map( a => p_1(6)(24), b => p_1(7)(24), cin => p_1(8)(24), cout => p_2(6)(25), s => p_2(2)(24)); 
fa_1_25_2: Full_Adder port map( a => p_1(6)(25), b => p_1(7)(25), cin => p_1(8)(25), cout => p_2(6)(26), s => p_2(2)(25)); 
fa_1_26_2: Full_Adder port map( a => p_1(6)(26), b => p_1(7)(26), cin => p_1(8)(26), cout => p_2(6)(27), s => p_2(2)(26)); 
fa_1_27_2: Full_Adder port map( a => p_1(6)(27), b => p_1(7)(27), cin => p_1(8)(27), cout => p_2(6)(28), s => p_2(2)(27)); 
fa_1_28_2: Full_Adder port map( a => p_1(6)(28), b => p_1(7)(28), cin => p_1(8)(28), cout => p_2(6)(29), s => p_2(2)(28)); 
fa_1_29_2: Full_Adder port map( a => p_1(6)(29), b => p_1(7)(29), cin => p_1(8)(29), cout => p_2(6)(30), s => p_2(2)(29)); 
fa_1_30_2: Full_Adder port map( a => p_1(6)(30), b => p_1(7)(30), cin => p_1(8)(30), cout => p_2(6)(31), s => p_2(2)(30)); 
fa_1_31_2: Full_Adder port map( a => p_1(6)(31), b => p_1(7)(31), cin => p_1(8)(31), cout => p_2(6)(32), s => p_2(2)(31)); 
fa_1_32_2: Full_Adder port map( a => p_1(6)(32), b => p_1(7)(32), cin => p_1(8)(32), cout => p_2(6)(33), s => p_2(2)(32)); 
fa_1_33_2: Full_Adder port map( a => p_1(6)(33), b => p_1(7)(33), cin => p_1(8)(33), cout => p_2(6)(34), s => p_2(2)(33)); 
fa_1_34_2: Full_Adder port map( a => p_1(6)(34), b => p_1(7)(34), cin => p_1(8)(34), cout => p_2(6)(35), s => p_2(2)(34)); 
fa_1_35_2: Full_Adder port map( a => p_1(6)(35), b => p_1(7)(35), cin => p_1(8)(35), cout => p_2(6)(36), s => p_2(2)(35)); 
fa_1_36_2: Full_Adder port map( a => p_1(6)(36), b => p_1(7)(36), cin => p_1(8)(36), cout => p_2(6)(37), s => p_2(2)(36)); 
fa_1_37_2: Full_Adder port map( a => p_1(6)(37), b => p_1(7)(37), cin => p_1(8)(37), cout => p_2(6)(38), s => p_2(2)(37)); 
fa_1_38_2: Full_Adder port map( a => p_1(6)(38), b => p_1(7)(38), cin => p_1(8)(38), cout => p_2(6)(39), s => p_2(2)(38)); 
fa_1_39_2: Full_Adder port map( a => p_1(6)(39), b => p_1(7)(39), cin => p_1(8)(39), cout => p_2(6)(40), s => p_2(2)(39)); 
fa_1_40_2: Full_Adder port map( a => p_1(6)(40), b => p_1(7)(40), cin => p_1(8)(40), cout => p_2(6)(41), s => p_2(2)(40)); 
fa_1_41_2: Full_Adder port map( a => p_1(6)(41), b => p_1(7)(41), cin => p_1(8)(41), cout => p_2(6)(42), s => p_2(2)(41)); 
fa_1_42_2: Full_Adder port map( a => p_1(6)(42), b => p_1(7)(42), cin => p_1(8)(42), cout => p_2(6)(43), s => p_2(2)(42)); 
fa_1_43_2: Full_Adder port map( a => p_1(6)(43), b => p_1(7)(43), cin => p_1(8)(43), cout => p_2(6)(44), s => p_2(2)(43)); 
fa_1_45_2: Full_Adder port map( a => p_1(6)(45), b => p_1(7)(45), cin => p_1(8)(45), cout => p_2(6)(46), s => p_2(2)(45)); 
p_2(2)(47) <= p_1(6)(47); 
p_2(3)(48) <= p_1(6)(48); 
p_2(4)(49) <= p_1(6)(49); 
p_2(5)(50) <= p_1(6)(50); 
p_2(6)(51) <= p_1(6)(51); 
p_2(6)(52) <= p_1(6)(52); 
p_2(6)(53) <= p_1(6)(53); 
p_2(6)(54) <= p_1(6)(54); 
p_2(7)(12) <= p_1(7)(12); 
p_2(7)(14) <= p_1(7)(14); 
p_2(7)(15) <= p_1(7)(15); 
p_2(6)(16) <= p_1(7)(16); 
p_2(6)(17) <= p_1(7)(17); 
p_2(4)(18) <= p_1(7)(18); 
p_2(4)(19) <= p_1(7)(19); 
p_2(3)(47) <= p_1(7)(47); 
p_2(4)(48) <= p_1(7)(48); 
p_2(5)(49) <= p_1(7)(49); 
p_2(6)(50) <= p_1(7)(50); 
p_2(7)(51) <= p_1(7)(51); 
p_2(7)(52) <= p_1(7)(52); 
p_2(8)(14) <= p_1(8)(14); 
p_2(7)(16) <= p_1(8)(16); 
p_2(7)(17) <= p_1(8)(17); 
p_2(5)(18) <= p_1(8)(18); 
p_2(5)(19) <= p_1(8)(19); 
p_2(3)(20) <= p_1(8)(20); 
p_2(3)(21) <= p_1(8)(21); 
fa_1_22_2: Full_Adder port map( a => p_1(8)(22), b => p_1(9)(22), cin => p_1(10)(22), cout => p_2(5)(23), s => p_2(3)(22)); 
fa_1_23_2: Full_Adder port map( a => p_1(8)(23), b => p_1(9)(23), cin => p_1(10)(23), cout => p_2(5)(24), s => p_2(3)(23)); 
fa_1_44_2: Full_Adder port map( a => p_1(8)(44), b => p_1(9)(44), cin => p_1(10)(44), cout => p_2(5)(45), s => p_2(3)(44)); 
p_2(3)(46) <= p_1(8)(46); 
p_2(4)(47) <= p_1(8)(47); 
p_2(5)(48) <= p_1(8)(48); 
p_2(6)(49) <= p_1(8)(49); 
p_2(7)(50) <= p_1(8)(50); 
p_2(8)(16) <= p_1(9)(16); 
p_2(6)(18) <= p_1(9)(18); 
p_2(6)(19) <= p_1(9)(19); 
p_2(4)(20) <= p_1(9)(20); 
p_2(4)(21) <= p_1(9)(21); 
fa_1_24_3: Full_Adder port map( a => p_1(9)(24), b => p_1(10)(24), cin => p_1(11)(24), cout => p_2(5)(25), s => p_2(3)(24)); 
fa_1_25_3: Full_Adder port map( a => p_1(9)(25), b => p_1(10)(25), cin => p_1(11)(25), cout => p_2(5)(26), s => p_2(3)(25)); 
fa_1_26_3: Full_Adder port map( a => p_1(9)(26), b => p_1(10)(26), cin => p_1(11)(26), cout => p_2(5)(27), s => p_2(3)(26)); 
fa_1_27_3: Full_Adder port map( a => p_1(9)(27), b => p_1(10)(27), cin => p_1(11)(27), cout => p_2(5)(28), s => p_2(3)(27)); 
fa_1_28_3: Full_Adder port map( a => p_1(9)(28), b => p_1(10)(28), cin => p_1(11)(28), cout => p_2(5)(29), s => p_2(3)(28)); 
fa_1_29_3: Full_Adder port map( a => p_1(9)(29), b => p_1(10)(29), cin => p_1(11)(29), cout => p_2(5)(30), s => p_2(3)(29)); 
fa_1_30_3: Full_Adder port map( a => p_1(9)(30), b => p_1(10)(30), cin => p_1(11)(30), cout => p_2(5)(31), s => p_2(3)(30)); 
fa_1_31_3: Full_Adder port map( a => p_1(9)(31), b => p_1(10)(31), cin => p_1(11)(31), cout => p_2(5)(32), s => p_2(3)(31)); 
fa_1_32_3: Full_Adder port map( a => p_1(9)(32), b => p_1(10)(32), cin => p_1(11)(32), cout => p_2(5)(33), s => p_2(3)(32)); 
fa_1_33_3: Full_Adder port map( a => p_1(9)(33), b => p_1(10)(33), cin => p_1(11)(33), cout => p_2(5)(34), s => p_2(3)(33)); 
fa_1_34_3: Full_Adder port map( a => p_1(9)(34), b => p_1(10)(34), cin => p_1(11)(34), cout => p_2(5)(35), s => p_2(3)(34)); 
fa_1_35_3: Full_Adder port map( a => p_1(9)(35), b => p_1(10)(35), cin => p_1(11)(35), cout => p_2(5)(36), s => p_2(3)(35)); 
fa_1_36_3: Full_Adder port map( a => p_1(9)(36), b => p_1(10)(36), cin => p_1(11)(36), cout => p_2(5)(37), s => p_2(3)(36)); 
fa_1_37_3: Full_Adder port map( a => p_1(9)(37), b => p_1(10)(37), cin => p_1(11)(37), cout => p_2(5)(38), s => p_2(3)(37)); 
fa_1_38_3: Full_Adder port map( a => p_1(9)(38), b => p_1(10)(38), cin => p_1(11)(38), cout => p_2(5)(39), s => p_2(3)(38)); 
fa_1_39_3: Full_Adder port map( a => p_1(9)(39), b => p_1(10)(39), cin => p_1(11)(39), cout => p_2(5)(40), s => p_2(3)(39)); 
fa_1_40_3: Full_Adder port map( a => p_1(9)(40), b => p_1(10)(40), cin => p_1(11)(40), cout => p_2(5)(41), s => p_2(3)(40)); 
fa_1_41_3: Full_Adder port map( a => p_1(9)(41), b => p_1(10)(41), cin => p_1(11)(41), cout => p_2(5)(42), s => p_2(3)(41)); 
fa_1_42_3: Full_Adder port map( a => p_1(9)(42), b => p_1(10)(42), cin => p_1(11)(42), cout => p_2(5)(43), s => p_2(3)(42)); 
fa_1_43_3: Full_Adder port map( a => p_1(9)(43), b => p_1(10)(43), cin => p_1(11)(43), cout => p_2(5)(44), s => p_2(3)(43)); 
p_2(3)(45) <= p_1(9)(45); 
p_2(4)(46) <= p_1(9)(46); 
p_2(5)(47) <= p_1(9)(47); 
p_2(6)(48) <= p_1(9)(48); 
p_2(7)(18) <= p_1(10)(18); 
p_2(5)(20) <= p_1(10)(20); 
p_2(5)(21) <= p_1(10)(21); 
p_2(4)(45) <= p_1(10)(45); 
p_2(5)(46) <= p_1(10)(46); 
p_2(6)(20) <= p_1(11)(20); 
p_2(4)(22) <= p_1(11)(22); 
p_2(4)(23) <= p_1(11)(23); 
p_2(4)(44) <= p_1(11)(44); 
p_2(5)(22) <= p_1(12)(22); 
p_2(4)(24) <= p_1(12)(24); 
p_2(4)(25) <= p_1(12)(25); 
p_2(4)(26) <= p_1(12)(26); 
p_2(4)(27) <= p_1(12)(27); 
p_2(4)(28) <= p_1(12)(28); 
p_2(4)(29) <= p_1(12)(29); 
p_2(4)(30) <= p_1(12)(30); 
p_2(4)(31) <= p_1(12)(31); 
p_2(4)(32) <= p_1(12)(32); 
p_2(4)(33) <= p_1(12)(33); 
p_2(4)(34) <= p_1(12)(34); 
p_2(4)(35) <= p_1(12)(35); 
p_2(4)(36) <= p_1(12)(36); 
p_2(4)(37) <= p_1(12)(37); 
p_2(4)(38) <= p_1(12)(38); 
p_2(4)(39) <= p_1(12)(39); 
p_2(4)(40) <= p_1(12)(40); 
p_2(4)(41) <= p_1(12)(41); 
p_2(4)(42) <= p_1(12)(42); 
p_2(4)(43) <= p_1(12)(43); 
p_3(0)(0) <= p_2(0)(0); 
p_3(0)(1) <= p_2(0)(1); 
p_3(0)(2) <= p_2(0)(2); 
p_3(0)(3) <= p_2(0)(3); 
p_3(0)(4) <= p_2(0)(4); 
p_3(0)(5) <= p_2(0)(5); 
p_3(0)(6) <= p_2(0)(6); 
p_3(0)(7) <= p_2(0)(7); 
p_3(0)(8) <= p_2(0)(8); 
p_3(0)(9) <= p_2(0)(9); 
ha_2_10_0: Half_Adder port map( a => p_2(0)(10), b => p_2(1)(10), cout => p_3(5)(11), s => p_3(0)(10)); 
ha_2_11_0: Half_Adder port map( a => p_2(0)(11), b => p_2(1)(11), cout => p_3(5)(12), s => p_3(0)(11)); 
ha_2_12_0: Half_Adder port map( a => p_2(0)(12), b => p_2(1)(12), cout => p_3(5)(13), s => p_3(0)(12)); 
ha_2_13_0: Half_Adder port map( a => p_2(0)(13), b => p_2(1)(13), cout => p_3(5)(14), s => p_3(0)(13)); 
ha_2_14_0: Half_Adder port map( a => p_2(0)(14), b => p_2(1)(14), cout => p_3(5)(15), s => p_3(0)(14)); 
ha_2_15_0: Half_Adder port map( a => p_2(0)(15), b => p_2(1)(15), cout => p_3(5)(16), s => p_3(0)(15)); 
fa_2_16_0: Full_Adder port map( a => p_2(0)(16), b => p_2(1)(16), cin => p_2(2)(16), cout => p_3(5)(17), s => p_3(0)(16)); 
fa_2_17_0: Full_Adder port map( a => p_2(0)(17), b => p_2(1)(17), cin => p_2(2)(17), cout => p_3(5)(18), s => p_3(0)(17)); 
fa_2_18_0: Full_Adder port map( a => p_2(0)(18), b => p_2(1)(18), cin => p_2(2)(18), cout => p_3(5)(19), s => p_3(0)(18)); 
fa_2_19_0: Full_Adder port map( a => p_2(0)(19), b => p_2(1)(19), cin => p_2(2)(19), cout => p_3(5)(20), s => p_3(0)(19)); 
fa_2_20_0: Full_Adder port map( a => p_2(0)(20), b => p_2(1)(20), cin => p_2(2)(20), cout => p_3(5)(21), s => p_3(0)(20)); 
fa_2_21_0: Full_Adder port map( a => p_2(0)(21), b => p_2(1)(21), cin => p_2(2)(21), cout => p_3(5)(22), s => p_3(0)(21)); 
fa_2_22_0: Full_Adder port map( a => p_2(0)(22), b => p_2(1)(22), cin => p_2(2)(22), cout => p_3(5)(23), s => p_3(0)(22)); 
fa_2_23_0: Full_Adder port map( a => p_2(0)(23), b => p_2(1)(23), cin => p_2(2)(23), cout => p_3(5)(24), s => p_3(0)(23)); 
fa_2_24_0: Full_Adder port map( a => p_2(0)(24), b => p_2(1)(24), cin => p_2(2)(24), cout => p_3(5)(25), s => p_3(0)(24)); 
fa_2_25_0: Full_Adder port map( a => p_2(0)(25), b => p_2(1)(25), cin => p_2(2)(25), cout => p_3(5)(26), s => p_3(0)(25)); 
fa_2_26_0: Full_Adder port map( a => p_2(0)(26), b => p_2(1)(26), cin => p_2(2)(26), cout => p_3(5)(27), s => p_3(0)(26)); 
fa_2_27_0: Full_Adder port map( a => p_2(0)(27), b => p_2(1)(27), cin => p_2(2)(27), cout => p_3(5)(28), s => p_3(0)(27)); 
fa_2_28_0: Full_Adder port map( a => p_2(0)(28), b => p_2(1)(28), cin => p_2(2)(28), cout => p_3(5)(29), s => p_3(0)(28)); 
fa_2_29_0: Full_Adder port map( a => p_2(0)(29), b => p_2(1)(29), cin => p_2(2)(29), cout => p_3(5)(30), s => p_3(0)(29)); 
fa_2_30_0: Full_Adder port map( a => p_2(0)(30), b => p_2(1)(30), cin => p_2(2)(30), cout => p_3(5)(31), s => p_3(0)(30)); 
fa_2_31_0: Full_Adder port map( a => p_2(0)(31), b => p_2(1)(31), cin => p_2(2)(31), cout => p_3(5)(32), s => p_3(0)(31)); 
fa_2_32_0: Full_Adder port map( a => p_2(0)(32), b => p_2(1)(32), cin => p_2(2)(32), cout => p_3(5)(33), s => p_3(0)(32)); 
fa_2_33_0: Full_Adder port map( a => p_2(0)(33), b => p_2(1)(33), cin => p_2(2)(33), cout => p_3(5)(34), s => p_3(0)(33)); 
fa_2_34_0: Full_Adder port map( a => p_2(0)(34), b => p_2(1)(34), cin => p_2(2)(34), cout => p_3(5)(35), s => p_3(0)(34)); 
fa_2_35_0: Full_Adder port map( a => p_2(0)(35), b => p_2(1)(35), cin => p_2(2)(35), cout => p_3(5)(36), s => p_3(0)(35)); 
fa_2_36_0: Full_Adder port map( a => p_2(0)(36), b => p_2(1)(36), cin => p_2(2)(36), cout => p_3(5)(37), s => p_3(0)(36)); 
fa_2_37_0: Full_Adder port map( a => p_2(0)(37), b => p_2(1)(37), cin => p_2(2)(37), cout => p_3(5)(38), s => p_3(0)(37)); 
fa_2_38_0: Full_Adder port map( a => p_2(0)(38), b => p_2(1)(38), cin => p_2(2)(38), cout => p_3(5)(39), s => p_3(0)(38)); 
fa_2_39_0: Full_Adder port map( a => p_2(0)(39), b => p_2(1)(39), cin => p_2(2)(39), cout => p_3(5)(40), s => p_3(0)(39)); 
fa_2_40_0: Full_Adder port map( a => p_2(0)(40), b => p_2(1)(40), cin => p_2(2)(40), cout => p_3(5)(41), s => p_3(0)(40)); 
fa_2_41_0: Full_Adder port map( a => p_2(0)(41), b => p_2(1)(41), cin => p_2(2)(41), cout => p_3(5)(42), s => p_3(0)(41)); 
fa_2_42_0: Full_Adder port map( a => p_2(0)(42), b => p_2(1)(42), cin => p_2(2)(42), cout => p_3(5)(43), s => p_3(0)(42)); 
fa_2_43_0: Full_Adder port map( a => p_2(0)(43), b => p_2(1)(43), cin => p_2(2)(43), cout => p_3(5)(44), s => p_3(0)(43)); 
fa_2_44_0: Full_Adder port map( a => p_2(0)(44), b => p_2(1)(44), cin => p_2(2)(44), cout => p_3(5)(45), s => p_3(0)(44)); 
fa_2_45_0: Full_Adder port map( a => p_2(0)(45), b => p_2(1)(45), cin => p_2(2)(45), cout => p_3(5)(46), s => p_3(0)(45)); 
fa_2_46_0: Full_Adder port map( a => p_2(0)(46), b => p_2(1)(46), cin => p_2(2)(46), cout => p_3(5)(47), s => p_3(0)(46)); 
fa_2_47_0: Full_Adder port map( a => p_2(0)(47), b => p_2(1)(47), cin => p_2(2)(47), cout => p_3(5)(48), s => p_3(0)(47)); 
fa_2_48_0: Full_Adder port map( a => p_2(0)(48), b => p_2(1)(48), cin => p_2(2)(48), cout => p_3(5)(49), s => p_3(0)(48)); 
fa_2_49_0: Full_Adder port map( a => p_2(0)(49), b => p_2(1)(49), cin => p_2(2)(49), cout => p_3(5)(50), s => p_3(0)(49)); 
fa_2_50_0: Full_Adder port map( a => p_2(0)(50), b => p_2(1)(50), cin => p_2(2)(50), cout => p_3(5)(51), s => p_3(0)(50)); 
fa_2_51_0: Full_Adder port map( a => p_2(0)(51), b => p_2(1)(51), cin => p_2(2)(51), cout => p_3(5)(52), s => p_3(0)(51)); 
ha_2_52_0: Half_Adder port map( a => p_2(0)(52), b => p_2(1)(52), cout => p_3(5)(53), s => p_3(0)(52)); 
fa_2_53_0: Full_Adder port map( a => p_2(0)(53), b => p_2(1)(53), cin => p_2(2)(53), cout => p_3(5)(54), s => p_3(0)(53)); 
ha_2_54_0: Half_Adder port map( a => p_2(0)(54), b => p_2(1)(54), cout => p_3(5)(55), s => p_3(0)(54)); 
fa_2_55_0: Full_Adder port map( a => p_2(0)(55), b => p_2(1)(55), cin => p_2(2)(55), cout => p_3(5)(56), s => p_3(0)(55)); 
ha_2_56_0: Half_Adder port map( a => p_2(0)(56), b => p_2(1)(56), cout => p_3(5)(57), s => p_3(0)(56)); 
p_3(0)(57) <= p_2(0)(57); 
p_3(0)(58) <= p_2(0)(58); 
p_3(0)(59) <= p_2(0)(59); 
p_3(0)(60) <= p_2(0)(60); 
p_3(0)(61) <= p_2(0)(61); 
p_3(0)(62) <= p_2(0)(62); 
p_3(0)(63) <= p_2(0)(63); 
p_3(1)(0) <= p_2(1)(0); 
p_3(1)(2) <= p_2(1)(2); 
p_3(1)(3) <= p_2(1)(3); 
p_3(1)(4) <= p_2(1)(4); 
p_3(1)(5) <= p_2(1)(5); 
p_3(1)(6) <= p_2(1)(6); 
p_3(1)(7) <= p_2(1)(7); 
p_3(1)(8) <= p_2(1)(8); 
p_3(1)(9) <= p_2(1)(9); 
p_3(1)(57) <= p_2(1)(57); 
p_3(1)(58) <= p_2(1)(58); 
p_3(1)(59) <= p_2(1)(59); 
p_3(1)(60) <= p_2(1)(60); 
p_3(1)(61) <= p_2(1)(61); 
p_3(1)(62) <= p_2(1)(62); 
p_3(1)(63) <= p_2(1)(63); 
p_3(2)(2) <= p_2(2)(2); 
p_3(2)(4) <= p_2(2)(4); 
p_3(2)(5) <= p_2(2)(5); 
p_3(2)(6) <= p_2(2)(6); 
p_3(2)(7) <= p_2(2)(7); 
p_3(2)(8) <= p_2(2)(8); 
p_3(2)(9) <= p_2(2)(9); 
p_3(1)(10) <= p_2(2)(10); 
p_3(1)(11) <= p_2(2)(11); 
fa_2_12_0: Full_Adder port map( a => p_2(2)(12), b => p_2(3)(12), cin => p_2(4)(12), cout => p_3(4)(13), s => p_3(1)(12)); 
fa_2_13_0: Full_Adder port map( a => p_2(2)(13), b => p_2(3)(13), cin => p_2(4)(13), cout => p_3(4)(14), s => p_3(1)(13)); 
fa_2_14_0: Full_Adder port map( a => p_2(2)(14), b => p_2(3)(14), cin => p_2(4)(14), cout => p_3(4)(15), s => p_3(1)(14)); 
fa_2_15_0: Full_Adder port map( a => p_2(2)(15), b => p_2(3)(15), cin => p_2(4)(15), cout => p_3(4)(16), s => p_3(1)(15)); 
fa_2_52_0: Full_Adder port map( a => p_2(2)(52), b => p_2(3)(52), cin => p_2(4)(52), cout => p_3(4)(53), s => p_3(1)(52)); 
fa_2_54_0: Full_Adder port map( a => p_2(2)(54), b => p_2(3)(54), cin => p_2(4)(54), cout => p_3(4)(55), s => p_3(1)(54)); 
p_3(1)(56) <= p_2(2)(56); 
p_3(2)(57) <= p_2(2)(57); 
p_3(2)(58) <= p_2(2)(58); 
p_3(2)(59) <= p_2(2)(59); 
p_3(2)(60) <= p_2(2)(60); 
p_3(2)(61) <= p_2(2)(61); 
p_3(2)(62) <= p_2(2)(62); 
p_3(3)(4) <= p_2(3)(4); 
p_3(3)(6) <= p_2(3)(6); 
p_3(3)(7) <= p_2(3)(7); 
p_3(3)(8) <= p_2(3)(8); 
p_3(3)(9) <= p_2(3)(9); 
p_3(2)(10) <= p_2(3)(10); 
p_3(2)(11) <= p_2(3)(11); 
fa_2_16_1: Full_Adder port map( a => p_2(3)(16), b => p_2(4)(16), cin => p_2(5)(16), cout => p_3(4)(17), s => p_3(1)(16)); 
fa_2_17_1: Full_Adder port map( a => p_2(3)(17), b => p_2(4)(17), cin => p_2(5)(17), cout => p_3(4)(18), s => p_3(1)(17)); 
fa_2_18_1: Full_Adder port map( a => p_2(3)(18), b => p_2(4)(18), cin => p_2(5)(18), cout => p_3(4)(19), s => p_3(1)(18)); 
fa_2_19_1: Full_Adder port map( a => p_2(3)(19), b => p_2(4)(19), cin => p_2(5)(19), cout => p_3(4)(20), s => p_3(1)(19)); 
fa_2_20_1: Full_Adder port map( a => p_2(3)(20), b => p_2(4)(20), cin => p_2(5)(20), cout => p_3(4)(21), s => p_3(1)(20)); 
fa_2_21_1: Full_Adder port map( a => p_2(3)(21), b => p_2(4)(21), cin => p_2(5)(21), cout => p_3(4)(22), s => p_3(1)(21)); 
fa_2_22_1: Full_Adder port map( a => p_2(3)(22), b => p_2(4)(22), cin => p_2(5)(22), cout => p_3(4)(23), s => p_3(1)(22)); 
fa_2_23_1: Full_Adder port map( a => p_2(3)(23), b => p_2(4)(23), cin => p_2(5)(23), cout => p_3(4)(24), s => p_3(1)(23)); 
fa_2_24_1: Full_Adder port map( a => p_2(3)(24), b => p_2(4)(24), cin => p_2(5)(24), cout => p_3(4)(25), s => p_3(1)(24)); 
fa_2_25_1: Full_Adder port map( a => p_2(3)(25), b => p_2(4)(25), cin => p_2(5)(25), cout => p_3(4)(26), s => p_3(1)(25)); 
fa_2_26_1: Full_Adder port map( a => p_2(3)(26), b => p_2(4)(26), cin => p_2(5)(26), cout => p_3(4)(27), s => p_3(1)(26)); 
fa_2_27_1: Full_Adder port map( a => p_2(3)(27), b => p_2(4)(27), cin => p_2(5)(27), cout => p_3(4)(28), s => p_3(1)(27)); 
fa_2_28_1: Full_Adder port map( a => p_2(3)(28), b => p_2(4)(28), cin => p_2(5)(28), cout => p_3(4)(29), s => p_3(1)(28)); 
fa_2_29_1: Full_Adder port map( a => p_2(3)(29), b => p_2(4)(29), cin => p_2(5)(29), cout => p_3(4)(30), s => p_3(1)(29)); 
fa_2_30_1: Full_Adder port map( a => p_2(3)(30), b => p_2(4)(30), cin => p_2(5)(30), cout => p_3(4)(31), s => p_3(1)(30)); 
fa_2_31_1: Full_Adder port map( a => p_2(3)(31), b => p_2(4)(31), cin => p_2(5)(31), cout => p_3(4)(32), s => p_3(1)(31)); 
fa_2_32_1: Full_Adder port map( a => p_2(3)(32), b => p_2(4)(32), cin => p_2(5)(32), cout => p_3(4)(33), s => p_3(1)(32)); 
fa_2_33_1: Full_Adder port map( a => p_2(3)(33), b => p_2(4)(33), cin => p_2(5)(33), cout => p_3(4)(34), s => p_3(1)(33)); 
fa_2_34_1: Full_Adder port map( a => p_2(3)(34), b => p_2(4)(34), cin => p_2(5)(34), cout => p_3(4)(35), s => p_3(1)(34)); 
fa_2_35_1: Full_Adder port map( a => p_2(3)(35), b => p_2(4)(35), cin => p_2(5)(35), cout => p_3(4)(36), s => p_3(1)(35)); 
fa_2_36_1: Full_Adder port map( a => p_2(3)(36), b => p_2(4)(36), cin => p_2(5)(36), cout => p_3(4)(37), s => p_3(1)(36)); 
fa_2_37_1: Full_Adder port map( a => p_2(3)(37), b => p_2(4)(37), cin => p_2(5)(37), cout => p_3(4)(38), s => p_3(1)(37)); 
fa_2_38_1: Full_Adder port map( a => p_2(3)(38), b => p_2(4)(38), cin => p_2(5)(38), cout => p_3(4)(39), s => p_3(1)(38)); 
fa_2_39_1: Full_Adder port map( a => p_2(3)(39), b => p_2(4)(39), cin => p_2(5)(39), cout => p_3(4)(40), s => p_3(1)(39)); 
fa_2_40_1: Full_Adder port map( a => p_2(3)(40), b => p_2(4)(40), cin => p_2(5)(40), cout => p_3(4)(41), s => p_3(1)(40)); 
fa_2_41_1: Full_Adder port map( a => p_2(3)(41), b => p_2(4)(41), cin => p_2(5)(41), cout => p_3(4)(42), s => p_3(1)(41)); 
fa_2_42_1: Full_Adder port map( a => p_2(3)(42), b => p_2(4)(42), cin => p_2(5)(42), cout => p_3(4)(43), s => p_3(1)(42)); 
fa_2_43_1: Full_Adder port map( a => p_2(3)(43), b => p_2(4)(43), cin => p_2(5)(43), cout => p_3(4)(44), s => p_3(1)(43)); 
fa_2_44_1: Full_Adder port map( a => p_2(3)(44), b => p_2(4)(44), cin => p_2(5)(44), cout => p_3(4)(45), s => p_3(1)(44)); 
fa_2_45_1: Full_Adder port map( a => p_2(3)(45), b => p_2(4)(45), cin => p_2(5)(45), cout => p_3(4)(46), s => p_3(1)(45)); 
fa_2_46_1: Full_Adder port map( a => p_2(3)(46), b => p_2(4)(46), cin => p_2(5)(46), cout => p_3(4)(47), s => p_3(1)(46)); 
fa_2_47_1: Full_Adder port map( a => p_2(3)(47), b => p_2(4)(47), cin => p_2(5)(47), cout => p_3(4)(48), s => p_3(1)(47)); 
fa_2_48_1: Full_Adder port map( a => p_2(3)(48), b => p_2(4)(48), cin => p_2(5)(48), cout => p_3(4)(49), s => p_3(1)(48)); 
fa_2_49_1: Full_Adder port map( a => p_2(3)(49), b => p_2(4)(49), cin => p_2(5)(49), cout => p_3(4)(50), s => p_3(1)(49)); 
fa_2_50_1: Full_Adder port map( a => p_2(3)(50), b => p_2(4)(50), cin => p_2(5)(50), cout => p_3(4)(51), s => p_3(1)(50)); 
fa_2_51_1: Full_Adder port map( a => p_2(3)(51), b => p_2(4)(51), cin => p_2(5)(51), cout => p_3(4)(52), s => p_3(1)(51)); 
fa_2_53_1: Full_Adder port map( a => p_2(3)(53), b => p_2(4)(53), cin => p_2(5)(53), cout => p_3(4)(54), s => p_3(1)(53)); 
p_3(1)(55) <= p_2(3)(55); 
p_3(2)(56) <= p_2(3)(56); 
p_3(3)(57) <= p_2(3)(57); 
p_3(3)(58) <= p_2(3)(58); 
p_3(3)(59) <= p_2(3)(59); 
p_3(3)(60) <= p_2(3)(60); 
p_3(4)(6) <= p_2(4)(6); 
p_3(4)(8) <= p_2(4)(8); 
p_3(4)(9) <= p_2(4)(9); 
p_3(3)(10) <= p_2(4)(10); 
p_3(3)(11) <= p_2(4)(11); 
p_3(2)(55) <= p_2(4)(55); 
p_3(3)(56) <= p_2(4)(56); 
p_3(4)(57) <= p_2(4)(57); 
p_3(4)(58) <= p_2(4)(58); 
p_3(5)(8) <= p_2(5)(8); 
p_3(4)(10) <= p_2(5)(10); 
p_3(4)(11) <= p_2(5)(11); 
p_3(2)(12) <= p_2(5)(12); 
p_3(2)(13) <= p_2(5)(13); 
fa_2_14_1: Full_Adder port map( a => p_2(5)(14), b => p_2(6)(14), cin => p_2(7)(14), cout => p_3(3)(15), s => p_3(2)(14)); 
fa_2_15_1: Full_Adder port map( a => p_2(5)(15), b => p_2(6)(15), cin => p_2(7)(15), cout => p_3(3)(16), s => p_3(2)(15)); 
fa_2_52_1: Full_Adder port map( a => p_2(5)(52), b => p_2(6)(52), cin => p_2(7)(52), cout => p_3(3)(53), s => p_3(2)(52)); 
p_3(2)(54) <= p_2(5)(54); 
p_3(3)(55) <= p_2(5)(55); 
p_3(4)(56) <= p_2(5)(56); 
p_3(5)(10) <= p_2(6)(10); 
p_3(3)(12) <= p_2(6)(12); 
p_3(3)(13) <= p_2(6)(13); 
fa_2_16_2: Full_Adder port map( a => p_2(6)(16), b => p_2(7)(16), cin => p_2(8)(16), cout => p_3(3)(17), s => p_3(2)(16)); 
fa_2_17_2: Full_Adder port map( a => p_2(6)(17), b => p_2(7)(17), cin => p_2(8)(17), cout => p_3(3)(18), s => p_3(2)(17)); 
fa_2_18_2: Full_Adder port map( a => p_2(6)(18), b => p_2(7)(18), cin => p_2(8)(18), cout => p_3(3)(19), s => p_3(2)(18)); 
fa_2_19_2: Full_Adder port map( a => p_2(6)(19), b => p_2(7)(19), cin => p_2(8)(19), cout => p_3(3)(20), s => p_3(2)(19)); 
fa_2_20_2: Full_Adder port map( a => p_2(6)(20), b => p_2(7)(20), cin => p_2(8)(20), cout => p_3(3)(21), s => p_3(2)(20)); 
fa_2_21_2: Full_Adder port map( a => p_2(6)(21), b => p_2(7)(21), cin => p_2(8)(21), cout => p_3(3)(22), s => p_3(2)(21)); 
fa_2_22_2: Full_Adder port map( a => p_2(6)(22), b => p_2(7)(22), cin => p_2(8)(22), cout => p_3(3)(23), s => p_3(2)(22)); 
fa_2_23_2: Full_Adder port map( a => p_2(6)(23), b => p_2(7)(23), cin => p_2(8)(23), cout => p_3(3)(24), s => p_3(2)(23)); 
fa_2_24_2: Full_Adder port map( a => p_2(6)(24), b => p_2(7)(24), cin => p_2(8)(24), cout => p_3(3)(25), s => p_3(2)(24)); 
fa_2_25_2: Full_Adder port map( a => p_2(6)(25), b => p_2(7)(25), cin => p_2(8)(25), cout => p_3(3)(26), s => p_3(2)(25)); 
fa_2_26_2: Full_Adder port map( a => p_2(6)(26), b => p_2(7)(26), cin => p_2(8)(26), cout => p_3(3)(27), s => p_3(2)(26)); 
fa_2_27_2: Full_Adder port map( a => p_2(6)(27), b => p_2(7)(27), cin => p_2(8)(27), cout => p_3(3)(28), s => p_3(2)(27)); 
fa_2_28_2: Full_Adder port map( a => p_2(6)(28), b => p_2(7)(28), cin => p_2(8)(28), cout => p_3(3)(29), s => p_3(2)(28)); 
fa_2_29_2: Full_Adder port map( a => p_2(6)(29), b => p_2(7)(29), cin => p_2(8)(29), cout => p_3(3)(30), s => p_3(2)(29)); 
fa_2_30_2: Full_Adder port map( a => p_2(6)(30), b => p_2(7)(30), cin => p_2(8)(30), cout => p_3(3)(31), s => p_3(2)(30)); 
fa_2_31_2: Full_Adder port map( a => p_2(6)(31), b => p_2(7)(31), cin => p_2(8)(31), cout => p_3(3)(32), s => p_3(2)(31)); 
fa_2_32_2: Full_Adder port map( a => p_2(6)(32), b => p_2(7)(32), cin => p_2(8)(32), cout => p_3(3)(33), s => p_3(2)(32)); 
fa_2_33_2: Full_Adder port map( a => p_2(6)(33), b => p_2(7)(33), cin => p_2(8)(33), cout => p_3(3)(34), s => p_3(2)(33)); 
fa_2_34_2: Full_Adder port map( a => p_2(6)(34), b => p_2(7)(34), cin => p_2(8)(34), cout => p_3(3)(35), s => p_3(2)(34)); 
fa_2_35_2: Full_Adder port map( a => p_2(6)(35), b => p_2(7)(35), cin => p_2(8)(35), cout => p_3(3)(36), s => p_3(2)(35)); 
fa_2_36_2: Full_Adder port map( a => p_2(6)(36), b => p_2(7)(36), cin => p_2(8)(36), cout => p_3(3)(37), s => p_3(2)(36)); 
fa_2_37_2: Full_Adder port map( a => p_2(6)(37), b => p_2(7)(37), cin => p_2(8)(37), cout => p_3(3)(38), s => p_3(2)(37)); 
fa_2_38_2: Full_Adder port map( a => p_2(6)(38), b => p_2(7)(38), cin => p_2(8)(38), cout => p_3(3)(39), s => p_3(2)(38)); 
fa_2_39_2: Full_Adder port map( a => p_2(6)(39), b => p_2(7)(39), cin => p_2(8)(39), cout => p_3(3)(40), s => p_3(2)(39)); 
fa_2_40_2: Full_Adder port map( a => p_2(6)(40), b => p_2(7)(40), cin => p_2(8)(40), cout => p_3(3)(41), s => p_3(2)(40)); 
fa_2_41_2: Full_Adder port map( a => p_2(6)(41), b => p_2(7)(41), cin => p_2(8)(41), cout => p_3(3)(42), s => p_3(2)(41)); 
fa_2_42_2: Full_Adder port map( a => p_2(6)(42), b => p_2(7)(42), cin => p_2(8)(42), cout => p_3(3)(43), s => p_3(2)(42)); 
fa_2_43_2: Full_Adder port map( a => p_2(6)(43), b => p_2(7)(43), cin => p_2(8)(43), cout => p_3(3)(44), s => p_3(2)(43)); 
fa_2_44_2: Full_Adder port map( a => p_2(6)(44), b => p_2(7)(44), cin => p_2(8)(44), cout => p_3(3)(45), s => p_3(2)(44)); 
fa_2_45_2: Full_Adder port map( a => p_2(6)(45), b => p_2(7)(45), cin => p_2(8)(45), cout => p_3(3)(46), s => p_3(2)(45)); 
fa_2_46_2: Full_Adder port map( a => p_2(6)(46), b => p_2(7)(46), cin => p_2(8)(46), cout => p_3(3)(47), s => p_3(2)(46)); 
fa_2_47_2: Full_Adder port map( a => p_2(6)(47), b => p_2(7)(47), cin => p_2(8)(47), cout => p_3(3)(48), s => p_3(2)(47)); 
fa_2_48_2: Full_Adder port map( a => p_2(6)(48), b => p_2(7)(48), cin => p_2(8)(48), cout => p_3(3)(49), s => p_3(2)(48)); 
fa_2_49_2: Full_Adder port map( a => p_2(6)(49), b => p_2(7)(49), cin => p_2(8)(49), cout => p_3(3)(50), s => p_3(2)(49)); 
fa_2_50_2: Full_Adder port map( a => p_2(6)(50), b => p_2(7)(50), cin => p_2(8)(50), cout => p_3(3)(51), s => p_3(2)(50)); 
fa_2_51_2: Full_Adder port map( a => p_2(6)(51), b => p_2(7)(51), cin => p_2(8)(51), cout => p_3(3)(52), s => p_3(2)(51)); 
p_3(2)(53) <= p_2(6)(53); 
p_3(3)(54) <= p_2(6)(54); 
p_3(4)(12) <= p_2(7)(12); 
p_3(3)(14) <= p_2(8)(14); 
p_4(0)(0) <= p_3(0)(0); 
p_4(0)(1) <= p_3(0)(1); 
p_4(0)(2) <= p_3(0)(2); 
p_4(0)(3) <= p_3(0)(3); 
p_4(0)(4) <= p_3(0)(4); 
p_4(0)(5) <= p_3(0)(5); 
ha_3_6_0: Half_Adder port map( a => p_3(0)(6), b => p_3(1)(6), cout => p_4(3)(7), s => p_4(0)(6)); 
ha_3_7_0: Half_Adder port map( a => p_3(0)(7), b => p_3(1)(7), cout => p_4(3)(8), s => p_4(0)(7)); 
ha_3_8_0: Half_Adder port map( a => p_3(0)(8), b => p_3(1)(8), cout => p_4(3)(9), s => p_4(0)(8)); 
ha_3_9_0: Half_Adder port map( a => p_3(0)(9), b => p_3(1)(9), cout => p_4(3)(10), s => p_4(0)(9)); 
fa_3_10_0: Full_Adder port map( a => p_3(0)(10), b => p_3(1)(10), cin => p_3(2)(10), cout => p_4(3)(11), s => p_4(0)(10)); 
fa_3_11_0: Full_Adder port map( a => p_3(0)(11), b => p_3(1)(11), cin => p_3(2)(11), cout => p_4(3)(12), s => p_4(0)(11)); 
fa_3_12_0: Full_Adder port map( a => p_3(0)(12), b => p_3(1)(12), cin => p_3(2)(12), cout => p_4(3)(13), s => p_4(0)(12)); 
fa_3_13_0: Full_Adder port map( a => p_3(0)(13), b => p_3(1)(13), cin => p_3(2)(13), cout => p_4(3)(14), s => p_4(0)(13)); 
fa_3_14_0: Full_Adder port map( a => p_3(0)(14), b => p_3(1)(14), cin => p_3(2)(14), cout => p_4(3)(15), s => p_4(0)(14)); 
fa_3_15_0: Full_Adder port map( a => p_3(0)(15), b => p_3(1)(15), cin => p_3(2)(15), cout => p_4(3)(16), s => p_4(0)(15)); 
fa_3_16_0: Full_Adder port map( a => p_3(0)(16), b => p_3(1)(16), cin => p_3(2)(16), cout => p_4(3)(17), s => p_4(0)(16)); 
fa_3_17_0: Full_Adder port map( a => p_3(0)(17), b => p_3(1)(17), cin => p_3(2)(17), cout => p_4(3)(18), s => p_4(0)(17)); 
fa_3_18_0: Full_Adder port map( a => p_3(0)(18), b => p_3(1)(18), cin => p_3(2)(18), cout => p_4(3)(19), s => p_4(0)(18)); 
fa_3_19_0: Full_Adder port map( a => p_3(0)(19), b => p_3(1)(19), cin => p_3(2)(19), cout => p_4(3)(20), s => p_4(0)(19)); 
fa_3_20_0: Full_Adder port map( a => p_3(0)(20), b => p_3(1)(20), cin => p_3(2)(20), cout => p_4(3)(21), s => p_4(0)(20)); 
fa_3_21_0: Full_Adder port map( a => p_3(0)(21), b => p_3(1)(21), cin => p_3(2)(21), cout => p_4(3)(22), s => p_4(0)(21)); 
fa_3_22_0: Full_Adder port map( a => p_3(0)(22), b => p_3(1)(22), cin => p_3(2)(22), cout => p_4(3)(23), s => p_4(0)(22)); 
fa_3_23_0: Full_Adder port map( a => p_3(0)(23), b => p_3(1)(23), cin => p_3(2)(23), cout => p_4(3)(24), s => p_4(0)(23)); 
fa_3_24_0: Full_Adder port map( a => p_3(0)(24), b => p_3(1)(24), cin => p_3(2)(24), cout => p_4(3)(25), s => p_4(0)(24)); 
fa_3_25_0: Full_Adder port map( a => p_3(0)(25), b => p_3(1)(25), cin => p_3(2)(25), cout => p_4(3)(26), s => p_4(0)(25)); 
fa_3_26_0: Full_Adder port map( a => p_3(0)(26), b => p_3(1)(26), cin => p_3(2)(26), cout => p_4(3)(27), s => p_4(0)(26)); 
fa_3_27_0: Full_Adder port map( a => p_3(0)(27), b => p_3(1)(27), cin => p_3(2)(27), cout => p_4(3)(28), s => p_4(0)(27)); 
fa_3_28_0: Full_Adder port map( a => p_3(0)(28), b => p_3(1)(28), cin => p_3(2)(28), cout => p_4(3)(29), s => p_4(0)(28)); 
fa_3_29_0: Full_Adder port map( a => p_3(0)(29), b => p_3(1)(29), cin => p_3(2)(29), cout => p_4(3)(30), s => p_4(0)(29)); 
fa_3_30_0: Full_Adder port map( a => p_3(0)(30), b => p_3(1)(30), cin => p_3(2)(30), cout => p_4(3)(31), s => p_4(0)(30)); 
fa_3_31_0: Full_Adder port map( a => p_3(0)(31), b => p_3(1)(31), cin => p_3(2)(31), cout => p_4(3)(32), s => p_4(0)(31)); 
fa_3_32_0: Full_Adder port map( a => p_3(0)(32), b => p_3(1)(32), cin => p_3(2)(32), cout => p_4(3)(33), s => p_4(0)(32)); 
fa_3_33_0: Full_Adder port map( a => p_3(0)(33), b => p_3(1)(33), cin => p_3(2)(33), cout => p_4(3)(34), s => p_4(0)(33)); 
fa_3_34_0: Full_Adder port map( a => p_3(0)(34), b => p_3(1)(34), cin => p_3(2)(34), cout => p_4(3)(35), s => p_4(0)(34)); 
fa_3_35_0: Full_Adder port map( a => p_3(0)(35), b => p_3(1)(35), cin => p_3(2)(35), cout => p_4(3)(36), s => p_4(0)(35)); 
fa_3_36_0: Full_Adder port map( a => p_3(0)(36), b => p_3(1)(36), cin => p_3(2)(36), cout => p_4(3)(37), s => p_4(0)(36)); 
fa_3_37_0: Full_Adder port map( a => p_3(0)(37), b => p_3(1)(37), cin => p_3(2)(37), cout => p_4(3)(38), s => p_4(0)(37)); 
fa_3_38_0: Full_Adder port map( a => p_3(0)(38), b => p_3(1)(38), cin => p_3(2)(38), cout => p_4(3)(39), s => p_4(0)(38)); 
fa_3_39_0: Full_Adder port map( a => p_3(0)(39), b => p_3(1)(39), cin => p_3(2)(39), cout => p_4(3)(40), s => p_4(0)(39)); 
fa_3_40_0: Full_Adder port map( a => p_3(0)(40), b => p_3(1)(40), cin => p_3(2)(40), cout => p_4(3)(41), s => p_4(0)(40)); 
fa_3_41_0: Full_Adder port map( a => p_3(0)(41), b => p_3(1)(41), cin => p_3(2)(41), cout => p_4(3)(42), s => p_4(0)(41)); 
fa_3_42_0: Full_Adder port map( a => p_3(0)(42), b => p_3(1)(42), cin => p_3(2)(42), cout => p_4(3)(43), s => p_4(0)(42)); 
fa_3_43_0: Full_Adder port map( a => p_3(0)(43), b => p_3(1)(43), cin => p_3(2)(43), cout => p_4(3)(44), s => p_4(0)(43)); 
fa_3_44_0: Full_Adder port map( a => p_3(0)(44), b => p_3(1)(44), cin => p_3(2)(44), cout => p_4(3)(45), s => p_4(0)(44)); 
fa_3_45_0: Full_Adder port map( a => p_3(0)(45), b => p_3(1)(45), cin => p_3(2)(45), cout => p_4(3)(46), s => p_4(0)(45)); 
fa_3_46_0: Full_Adder port map( a => p_3(0)(46), b => p_3(1)(46), cin => p_3(2)(46), cout => p_4(3)(47), s => p_4(0)(46)); 
fa_3_47_0: Full_Adder port map( a => p_3(0)(47), b => p_3(1)(47), cin => p_3(2)(47), cout => p_4(3)(48), s => p_4(0)(47)); 
fa_3_48_0: Full_Adder port map( a => p_3(0)(48), b => p_3(1)(48), cin => p_3(2)(48), cout => p_4(3)(49), s => p_4(0)(48)); 
fa_3_49_0: Full_Adder port map( a => p_3(0)(49), b => p_3(1)(49), cin => p_3(2)(49), cout => p_4(3)(50), s => p_4(0)(49)); 
fa_3_50_0: Full_Adder port map( a => p_3(0)(50), b => p_3(1)(50), cin => p_3(2)(50), cout => p_4(3)(51), s => p_4(0)(50)); 
fa_3_51_0: Full_Adder port map( a => p_3(0)(51), b => p_3(1)(51), cin => p_3(2)(51), cout => p_4(3)(52), s => p_4(0)(51)); 
fa_3_52_0: Full_Adder port map( a => p_3(0)(52), b => p_3(1)(52), cin => p_3(2)(52), cout => p_4(3)(53), s => p_4(0)(52)); 
fa_3_53_0: Full_Adder port map( a => p_3(0)(53), b => p_3(1)(53), cin => p_3(2)(53), cout => p_4(3)(54), s => p_4(0)(53)); 
fa_3_54_0: Full_Adder port map( a => p_3(0)(54), b => p_3(1)(54), cin => p_3(2)(54), cout => p_4(3)(55), s => p_4(0)(54)); 
fa_3_55_0: Full_Adder port map( a => p_3(0)(55), b => p_3(1)(55), cin => p_3(2)(55), cout => p_4(3)(56), s => p_4(0)(55)); 
fa_3_56_0: Full_Adder port map( a => p_3(0)(56), b => p_3(1)(56), cin => p_3(2)(56), cout => p_4(3)(57), s => p_4(0)(56)); 
fa_3_57_0: Full_Adder port map( a => p_3(0)(57), b => p_3(1)(57), cin => p_3(2)(57), cout => p_4(3)(58), s => p_4(0)(57)); 
ha_3_58_0: Half_Adder port map( a => p_3(0)(58), b => p_3(1)(58), cout => p_4(3)(59), s => p_4(0)(58)); 
fa_3_59_0: Full_Adder port map( a => p_3(0)(59), b => p_3(1)(59), cin => p_3(2)(59), cout => p_4(3)(60), s => p_4(0)(59)); 
ha_3_60_0: Half_Adder port map( a => p_3(0)(60), b => p_3(1)(60), cout => p_4(3)(61), s => p_4(0)(60)); 
p_4(0)(61) <= p_3(0)(61); 
p_4(0)(62) <= p_3(0)(62); 
p_4(0)(63) <= p_3(0)(63); 
p_4(1)(0) <= p_3(1)(0); 
p_4(1)(2) <= p_3(1)(2); 
p_4(1)(3) <= p_3(1)(3); 
p_4(1)(4) <= p_3(1)(4); 
p_4(1)(5) <= p_3(1)(5); 
p_4(1)(61) <= p_3(1)(61); 
p_4(1)(62) <= p_3(1)(62); 
p_4(1)(63) <= p_3(1)(63); 
p_4(2)(2) <= p_3(2)(2); 
p_4(2)(4) <= p_3(2)(4); 
p_4(2)(5) <= p_3(2)(5); 
p_4(1)(6) <= p_3(2)(6); 
p_4(1)(7) <= p_3(2)(7); 
fa_3_8_0: Full_Adder port map( a => p_3(2)(8), b => p_3(3)(8), cin => p_3(4)(8), cout => p_4(2)(9), s => p_4(1)(8)); 
fa_3_9_0: Full_Adder port map( a => p_3(2)(9), b => p_3(3)(9), cin => p_3(4)(9), cout => p_4(2)(10), s => p_4(1)(9)); 
fa_3_58_0: Full_Adder port map( a => p_3(2)(58), b => p_3(3)(58), cin => p_3(4)(58), cout => p_4(2)(59), s => p_4(1)(58)); 
p_4(1)(60) <= p_3(2)(60); 
p_4(2)(61) <= p_3(2)(61); 
p_4(2)(62) <= p_3(2)(62); 
p_4(3)(4) <= p_3(3)(4); 
p_4(2)(6) <= p_3(3)(6); 
p_4(2)(7) <= p_3(3)(7); 
fa_3_10_1: Full_Adder port map( a => p_3(3)(10), b => p_3(4)(10), cin => p_3(5)(10), cout => p_4(2)(11), s => p_4(1)(10)); 
fa_3_11_1: Full_Adder port map( a => p_3(3)(11), b => p_3(4)(11), cin => p_3(5)(11), cout => p_4(2)(12), s => p_4(1)(11)); 
fa_3_12_1: Full_Adder port map( a => p_3(3)(12), b => p_3(4)(12), cin => p_3(5)(12), cout => p_4(2)(13), s => p_4(1)(12)); 
fa_3_13_1: Full_Adder port map( a => p_3(3)(13), b => p_3(4)(13), cin => p_3(5)(13), cout => p_4(2)(14), s => p_4(1)(13)); 
fa_3_14_1: Full_Adder port map( a => p_3(3)(14), b => p_3(4)(14), cin => p_3(5)(14), cout => p_4(2)(15), s => p_4(1)(14)); 
fa_3_15_1: Full_Adder port map( a => p_3(3)(15), b => p_3(4)(15), cin => p_3(5)(15), cout => p_4(2)(16), s => p_4(1)(15)); 
fa_3_16_1: Full_Adder port map( a => p_3(3)(16), b => p_3(4)(16), cin => p_3(5)(16), cout => p_4(2)(17), s => p_4(1)(16)); 
fa_3_17_1: Full_Adder port map( a => p_3(3)(17), b => p_3(4)(17), cin => p_3(5)(17), cout => p_4(2)(18), s => p_4(1)(17)); 
fa_3_18_1: Full_Adder port map( a => p_3(3)(18), b => p_3(4)(18), cin => p_3(5)(18), cout => p_4(2)(19), s => p_4(1)(18)); 
fa_3_19_1: Full_Adder port map( a => p_3(3)(19), b => p_3(4)(19), cin => p_3(5)(19), cout => p_4(2)(20), s => p_4(1)(19)); 
fa_3_20_1: Full_Adder port map( a => p_3(3)(20), b => p_3(4)(20), cin => p_3(5)(20), cout => p_4(2)(21), s => p_4(1)(20)); 
fa_3_21_1: Full_Adder port map( a => p_3(3)(21), b => p_3(4)(21), cin => p_3(5)(21), cout => p_4(2)(22), s => p_4(1)(21)); 
fa_3_22_1: Full_Adder port map( a => p_3(3)(22), b => p_3(4)(22), cin => p_3(5)(22), cout => p_4(2)(23), s => p_4(1)(22)); 
fa_3_23_1: Full_Adder port map( a => p_3(3)(23), b => p_3(4)(23), cin => p_3(5)(23), cout => p_4(2)(24), s => p_4(1)(23)); 
fa_3_24_1: Full_Adder port map( a => p_3(3)(24), b => p_3(4)(24), cin => p_3(5)(24), cout => p_4(2)(25), s => p_4(1)(24)); 
fa_3_25_1: Full_Adder port map( a => p_3(3)(25), b => p_3(4)(25), cin => p_3(5)(25), cout => p_4(2)(26), s => p_4(1)(25)); 
fa_3_26_1: Full_Adder port map( a => p_3(3)(26), b => p_3(4)(26), cin => p_3(5)(26), cout => p_4(2)(27), s => p_4(1)(26)); 
fa_3_27_1: Full_Adder port map( a => p_3(3)(27), b => p_3(4)(27), cin => p_3(5)(27), cout => p_4(2)(28), s => p_4(1)(27)); 
fa_3_28_1: Full_Adder port map( a => p_3(3)(28), b => p_3(4)(28), cin => p_3(5)(28), cout => p_4(2)(29), s => p_4(1)(28)); 
fa_3_29_1: Full_Adder port map( a => p_3(3)(29), b => p_3(4)(29), cin => p_3(5)(29), cout => p_4(2)(30), s => p_4(1)(29)); 
fa_3_30_1: Full_Adder port map( a => p_3(3)(30), b => p_3(4)(30), cin => p_3(5)(30), cout => p_4(2)(31), s => p_4(1)(30)); 
fa_3_31_1: Full_Adder port map( a => p_3(3)(31), b => p_3(4)(31), cin => p_3(5)(31), cout => p_4(2)(32), s => p_4(1)(31)); 
fa_3_32_1: Full_Adder port map( a => p_3(3)(32), b => p_3(4)(32), cin => p_3(5)(32), cout => p_4(2)(33), s => p_4(1)(32)); 
fa_3_33_1: Full_Adder port map( a => p_3(3)(33), b => p_3(4)(33), cin => p_3(5)(33), cout => p_4(2)(34), s => p_4(1)(33)); 
fa_3_34_1: Full_Adder port map( a => p_3(3)(34), b => p_3(4)(34), cin => p_3(5)(34), cout => p_4(2)(35), s => p_4(1)(34)); 
fa_3_35_1: Full_Adder port map( a => p_3(3)(35), b => p_3(4)(35), cin => p_3(5)(35), cout => p_4(2)(36), s => p_4(1)(35)); 
fa_3_36_1: Full_Adder port map( a => p_3(3)(36), b => p_3(4)(36), cin => p_3(5)(36), cout => p_4(2)(37), s => p_4(1)(36)); 
fa_3_37_1: Full_Adder port map( a => p_3(3)(37), b => p_3(4)(37), cin => p_3(5)(37), cout => p_4(2)(38), s => p_4(1)(37)); 
fa_3_38_1: Full_Adder port map( a => p_3(3)(38), b => p_3(4)(38), cin => p_3(5)(38), cout => p_4(2)(39), s => p_4(1)(38)); 
fa_3_39_1: Full_Adder port map( a => p_3(3)(39), b => p_3(4)(39), cin => p_3(5)(39), cout => p_4(2)(40), s => p_4(1)(39)); 
fa_3_40_1: Full_Adder port map( a => p_3(3)(40), b => p_3(4)(40), cin => p_3(5)(40), cout => p_4(2)(41), s => p_4(1)(40)); 
fa_3_41_1: Full_Adder port map( a => p_3(3)(41), b => p_3(4)(41), cin => p_3(5)(41), cout => p_4(2)(42), s => p_4(1)(41)); 
fa_3_42_1: Full_Adder port map( a => p_3(3)(42), b => p_3(4)(42), cin => p_3(5)(42), cout => p_4(2)(43), s => p_4(1)(42)); 
fa_3_43_1: Full_Adder port map( a => p_3(3)(43), b => p_3(4)(43), cin => p_3(5)(43), cout => p_4(2)(44), s => p_4(1)(43)); 
fa_3_44_1: Full_Adder port map( a => p_3(3)(44), b => p_3(4)(44), cin => p_3(5)(44), cout => p_4(2)(45), s => p_4(1)(44)); 
fa_3_45_1: Full_Adder port map( a => p_3(3)(45), b => p_3(4)(45), cin => p_3(5)(45), cout => p_4(2)(46), s => p_4(1)(45)); 
fa_3_46_1: Full_Adder port map( a => p_3(3)(46), b => p_3(4)(46), cin => p_3(5)(46), cout => p_4(2)(47), s => p_4(1)(46)); 
fa_3_47_1: Full_Adder port map( a => p_3(3)(47), b => p_3(4)(47), cin => p_3(5)(47), cout => p_4(2)(48), s => p_4(1)(47)); 
fa_3_48_1: Full_Adder port map( a => p_3(3)(48), b => p_3(4)(48), cin => p_3(5)(48), cout => p_4(2)(49), s => p_4(1)(48)); 
fa_3_49_1: Full_Adder port map( a => p_3(3)(49), b => p_3(4)(49), cin => p_3(5)(49), cout => p_4(2)(50), s => p_4(1)(49)); 
fa_3_50_1: Full_Adder port map( a => p_3(3)(50), b => p_3(4)(50), cin => p_3(5)(50), cout => p_4(2)(51), s => p_4(1)(50)); 
fa_3_51_1: Full_Adder port map( a => p_3(3)(51), b => p_3(4)(51), cin => p_3(5)(51), cout => p_4(2)(52), s => p_4(1)(51)); 
fa_3_52_1: Full_Adder port map( a => p_3(3)(52), b => p_3(4)(52), cin => p_3(5)(52), cout => p_4(2)(53), s => p_4(1)(52)); 
fa_3_53_1: Full_Adder port map( a => p_3(3)(53), b => p_3(4)(53), cin => p_3(5)(53), cout => p_4(2)(54), s => p_4(1)(53)); 
fa_3_54_1: Full_Adder port map( a => p_3(3)(54), b => p_3(4)(54), cin => p_3(5)(54), cout => p_4(2)(55), s => p_4(1)(54)); 
fa_3_55_1: Full_Adder port map( a => p_3(3)(55), b => p_3(4)(55), cin => p_3(5)(55), cout => p_4(2)(56), s => p_4(1)(55)); 
fa_3_56_1: Full_Adder port map( a => p_3(3)(56), b => p_3(4)(56), cin => p_3(5)(56), cout => p_4(2)(57), s => p_4(1)(56)); 
fa_3_57_1: Full_Adder port map( a => p_3(3)(57), b => p_3(4)(57), cin => p_3(5)(57), cout => p_4(2)(58), s => p_4(1)(57)); 
p_4(1)(59) <= p_3(3)(59); 
p_4(2)(60) <= p_3(3)(60); 
p_4(3)(6) <= p_3(4)(6); 
p_4(2)(8) <= p_3(5)(8); 
p_5(0)(0) <= p_4(0)(0); 
p_5(0)(1) <= p_4(0)(1); 
p_5(0)(2) <= p_4(0)(2); 
p_5(0)(3) <= p_4(0)(3); 
ha_4_4_0: Half_Adder port map( a => p_4(0)(4), b => p_4(1)(4), cout => p_5(2)(5), s => p_5(0)(4)); 
ha_4_5_0: Half_Adder port map( a => p_4(0)(5), b => p_4(1)(5), cout => p_5(2)(6), s => p_5(0)(5)); 
fa_4_6_0: Full_Adder port map( a => p_4(0)(6), b => p_4(1)(6), cin => p_4(2)(6), cout => p_5(2)(7), s => p_5(0)(6)); 
fa_4_7_0: Full_Adder port map( a => p_4(0)(7), b => p_4(1)(7), cin => p_4(2)(7), cout => p_5(2)(8), s => p_5(0)(7)); 
fa_4_8_0: Full_Adder port map( a => p_4(0)(8), b => p_4(1)(8), cin => p_4(2)(8), cout => p_5(2)(9), s => p_5(0)(8)); 
fa_4_9_0: Full_Adder port map( a => p_4(0)(9), b => p_4(1)(9), cin => p_4(2)(9), cout => p_5(2)(10), s => p_5(0)(9)); 
fa_4_10_0: Full_Adder port map( a => p_4(0)(10), b => p_4(1)(10), cin => p_4(2)(10), cout => p_5(2)(11), s => p_5(0)(10)); 
fa_4_11_0: Full_Adder port map( a => p_4(0)(11), b => p_4(1)(11), cin => p_4(2)(11), cout => p_5(2)(12), s => p_5(0)(11)); 
fa_4_12_0: Full_Adder port map( a => p_4(0)(12), b => p_4(1)(12), cin => p_4(2)(12), cout => p_5(2)(13), s => p_5(0)(12)); 
fa_4_13_0: Full_Adder port map( a => p_4(0)(13), b => p_4(1)(13), cin => p_4(2)(13), cout => p_5(2)(14), s => p_5(0)(13)); 
fa_4_14_0: Full_Adder port map( a => p_4(0)(14), b => p_4(1)(14), cin => p_4(2)(14), cout => p_5(2)(15), s => p_5(0)(14)); 
fa_4_15_0: Full_Adder port map( a => p_4(0)(15), b => p_4(1)(15), cin => p_4(2)(15), cout => p_5(2)(16), s => p_5(0)(15)); 
fa_4_16_0: Full_Adder port map( a => p_4(0)(16), b => p_4(1)(16), cin => p_4(2)(16), cout => p_5(2)(17), s => p_5(0)(16)); 
fa_4_17_0: Full_Adder port map( a => p_4(0)(17), b => p_4(1)(17), cin => p_4(2)(17), cout => p_5(2)(18), s => p_5(0)(17)); 
fa_4_18_0: Full_Adder port map( a => p_4(0)(18), b => p_4(1)(18), cin => p_4(2)(18), cout => p_5(2)(19), s => p_5(0)(18)); 
fa_4_19_0: Full_Adder port map( a => p_4(0)(19), b => p_4(1)(19), cin => p_4(2)(19), cout => p_5(2)(20), s => p_5(0)(19)); 
fa_4_20_0: Full_Adder port map( a => p_4(0)(20), b => p_4(1)(20), cin => p_4(2)(20), cout => p_5(2)(21), s => p_5(0)(20)); 
fa_4_21_0: Full_Adder port map( a => p_4(0)(21), b => p_4(1)(21), cin => p_4(2)(21), cout => p_5(2)(22), s => p_5(0)(21)); 
fa_4_22_0: Full_Adder port map( a => p_4(0)(22), b => p_4(1)(22), cin => p_4(2)(22), cout => p_5(2)(23), s => p_5(0)(22)); 
fa_4_23_0: Full_Adder port map( a => p_4(0)(23), b => p_4(1)(23), cin => p_4(2)(23), cout => p_5(2)(24), s => p_5(0)(23)); 
fa_4_24_0: Full_Adder port map( a => p_4(0)(24), b => p_4(1)(24), cin => p_4(2)(24), cout => p_5(2)(25), s => p_5(0)(24)); 
fa_4_25_0: Full_Adder port map( a => p_4(0)(25), b => p_4(1)(25), cin => p_4(2)(25), cout => p_5(2)(26), s => p_5(0)(25)); 
fa_4_26_0: Full_Adder port map( a => p_4(0)(26), b => p_4(1)(26), cin => p_4(2)(26), cout => p_5(2)(27), s => p_5(0)(26)); 
fa_4_27_0: Full_Adder port map( a => p_4(0)(27), b => p_4(1)(27), cin => p_4(2)(27), cout => p_5(2)(28), s => p_5(0)(27)); 
fa_4_28_0: Full_Adder port map( a => p_4(0)(28), b => p_4(1)(28), cin => p_4(2)(28), cout => p_5(2)(29), s => p_5(0)(28)); 
fa_4_29_0: Full_Adder port map( a => p_4(0)(29), b => p_4(1)(29), cin => p_4(2)(29), cout => p_5(2)(30), s => p_5(0)(29)); 
fa_4_30_0: Full_Adder port map( a => p_4(0)(30), b => p_4(1)(30), cin => p_4(2)(30), cout => p_5(2)(31), s => p_5(0)(30)); 
fa_4_31_0: Full_Adder port map( a => p_4(0)(31), b => p_4(1)(31), cin => p_4(2)(31), cout => p_5(2)(32), s => p_5(0)(31)); 
fa_4_32_0: Full_Adder port map( a => p_4(0)(32), b => p_4(1)(32), cin => p_4(2)(32), cout => p_5(2)(33), s => p_5(0)(32)); 
fa_4_33_0: Full_Adder port map( a => p_4(0)(33), b => p_4(1)(33), cin => p_4(2)(33), cout => p_5(2)(34), s => p_5(0)(33)); 
fa_4_34_0: Full_Adder port map( a => p_4(0)(34), b => p_4(1)(34), cin => p_4(2)(34), cout => p_5(2)(35), s => p_5(0)(34)); 
fa_4_35_0: Full_Adder port map( a => p_4(0)(35), b => p_4(1)(35), cin => p_4(2)(35), cout => p_5(2)(36), s => p_5(0)(35)); 
fa_4_36_0: Full_Adder port map( a => p_4(0)(36), b => p_4(1)(36), cin => p_4(2)(36), cout => p_5(2)(37), s => p_5(0)(36)); 
fa_4_37_0: Full_Adder port map( a => p_4(0)(37), b => p_4(1)(37), cin => p_4(2)(37), cout => p_5(2)(38), s => p_5(0)(37)); 
fa_4_38_0: Full_Adder port map( a => p_4(0)(38), b => p_4(1)(38), cin => p_4(2)(38), cout => p_5(2)(39), s => p_5(0)(38)); 
fa_4_39_0: Full_Adder port map( a => p_4(0)(39), b => p_4(1)(39), cin => p_4(2)(39), cout => p_5(2)(40), s => p_5(0)(39)); 
fa_4_40_0: Full_Adder port map( a => p_4(0)(40), b => p_4(1)(40), cin => p_4(2)(40), cout => p_5(2)(41), s => p_5(0)(40)); 
fa_4_41_0: Full_Adder port map( a => p_4(0)(41), b => p_4(1)(41), cin => p_4(2)(41), cout => p_5(2)(42), s => p_5(0)(41)); 
fa_4_42_0: Full_Adder port map( a => p_4(0)(42), b => p_4(1)(42), cin => p_4(2)(42), cout => p_5(2)(43), s => p_5(0)(42)); 
fa_4_43_0: Full_Adder port map( a => p_4(0)(43), b => p_4(1)(43), cin => p_4(2)(43), cout => p_5(2)(44), s => p_5(0)(43)); 
fa_4_44_0: Full_Adder port map( a => p_4(0)(44), b => p_4(1)(44), cin => p_4(2)(44), cout => p_5(2)(45), s => p_5(0)(44)); 
fa_4_45_0: Full_Adder port map( a => p_4(0)(45), b => p_4(1)(45), cin => p_4(2)(45), cout => p_5(2)(46), s => p_5(0)(45)); 
fa_4_46_0: Full_Adder port map( a => p_4(0)(46), b => p_4(1)(46), cin => p_4(2)(46), cout => p_5(2)(47), s => p_5(0)(46)); 
fa_4_47_0: Full_Adder port map( a => p_4(0)(47), b => p_4(1)(47), cin => p_4(2)(47), cout => p_5(2)(48), s => p_5(0)(47)); 
fa_4_48_0: Full_Adder port map( a => p_4(0)(48), b => p_4(1)(48), cin => p_4(2)(48), cout => p_5(2)(49), s => p_5(0)(48)); 
fa_4_49_0: Full_Adder port map( a => p_4(0)(49), b => p_4(1)(49), cin => p_4(2)(49), cout => p_5(2)(50), s => p_5(0)(49)); 
fa_4_50_0: Full_Adder port map( a => p_4(0)(50), b => p_4(1)(50), cin => p_4(2)(50), cout => p_5(2)(51), s => p_5(0)(50)); 
fa_4_51_0: Full_Adder port map( a => p_4(0)(51), b => p_4(1)(51), cin => p_4(2)(51), cout => p_5(2)(52), s => p_5(0)(51)); 
fa_4_52_0: Full_Adder port map( a => p_4(0)(52), b => p_4(1)(52), cin => p_4(2)(52), cout => p_5(2)(53), s => p_5(0)(52)); 
fa_4_53_0: Full_Adder port map( a => p_4(0)(53), b => p_4(1)(53), cin => p_4(2)(53), cout => p_5(2)(54), s => p_5(0)(53)); 
fa_4_54_0: Full_Adder port map( a => p_4(0)(54), b => p_4(1)(54), cin => p_4(2)(54), cout => p_5(2)(55), s => p_5(0)(54)); 
fa_4_55_0: Full_Adder port map( a => p_4(0)(55), b => p_4(1)(55), cin => p_4(2)(55), cout => p_5(2)(56), s => p_5(0)(55)); 
fa_4_56_0: Full_Adder port map( a => p_4(0)(56), b => p_4(1)(56), cin => p_4(2)(56), cout => p_5(2)(57), s => p_5(0)(56)); 
fa_4_57_0: Full_Adder port map( a => p_4(0)(57), b => p_4(1)(57), cin => p_4(2)(57), cout => p_5(2)(58), s => p_5(0)(57)); 
fa_4_58_0: Full_Adder port map( a => p_4(0)(58), b => p_4(1)(58), cin => p_4(2)(58), cout => p_5(2)(59), s => p_5(0)(58)); 
fa_4_59_0: Full_Adder port map( a => p_4(0)(59), b => p_4(1)(59), cin => p_4(2)(59), cout => p_5(2)(60), s => p_5(0)(59)); 
fa_4_60_0: Full_Adder port map( a => p_4(0)(60), b => p_4(1)(60), cin => p_4(2)(60), cout => p_5(2)(61), s => p_5(0)(60)); 
fa_4_61_0: Full_Adder port map( a => p_4(0)(61), b => p_4(1)(61), cin => p_4(2)(61), cout => p_5(2)(62), s => p_5(0)(61)); 
ha_4_62_0: Half_Adder port map( a => p_4(0)(62), b => p_4(1)(62), cout => p_5(2)(63), s => p_5(0)(62)); 
p_5(0)(63) <= p_4(0)(63); 
p_5(1)(0) <= p_4(1)(0); 
p_5(1)(2) <= p_4(1)(2); 
p_5(1)(3) <= p_4(1)(3); 
p_5(1)(63) <= p_4(1)(63); 
p_5(2)(2) <= p_4(2)(2); 
p_5(1)(4) <= p_4(2)(4); 
p_5(1)(5) <= p_4(2)(5); 
p_5(1)(62) <= p_4(2)(62); 
p_5(2)(4) <= p_4(3)(4); 
p_5(1)(6) <= p_4(3)(6); 
p_5(1)(7) <= p_4(3)(7); 
p_5(1)(8) <= p_4(3)(8); 
p_5(1)(9) <= p_4(3)(9); 
p_5(1)(10) <= p_4(3)(10); 
p_5(1)(11) <= p_4(3)(11); 
p_5(1)(12) <= p_4(3)(12); 
p_5(1)(13) <= p_4(3)(13); 
p_5(1)(14) <= p_4(3)(14); 
p_5(1)(15) <= p_4(3)(15); 
p_5(1)(16) <= p_4(3)(16); 
p_5(1)(17) <= p_4(3)(17); 
p_5(1)(18) <= p_4(3)(18); 
p_5(1)(19) <= p_4(3)(19); 
p_5(1)(20) <= p_4(3)(20); 
p_5(1)(21) <= p_4(3)(21); 
p_5(1)(22) <= p_4(3)(22); 
p_5(1)(23) <= p_4(3)(23); 
p_5(1)(24) <= p_4(3)(24); 
p_5(1)(25) <= p_4(3)(25); 
p_5(1)(26) <= p_4(3)(26); 
p_5(1)(27) <= p_4(3)(27); 
p_5(1)(28) <= p_4(3)(28); 
p_5(1)(29) <= p_4(3)(29); 
p_5(1)(30) <= p_4(3)(30); 
p_5(1)(31) <= p_4(3)(31); 
p_5(1)(32) <= p_4(3)(32); 
p_5(1)(33) <= p_4(3)(33); 
p_5(1)(34) <= p_4(3)(34); 
p_5(1)(35) <= p_4(3)(35); 
p_5(1)(36) <= p_4(3)(36); 
p_5(1)(37) <= p_4(3)(37); 
p_5(1)(38) <= p_4(3)(38); 
p_5(1)(39) <= p_4(3)(39); 
p_5(1)(40) <= p_4(3)(40); 
p_5(1)(41) <= p_4(3)(41); 
p_5(1)(42) <= p_4(3)(42); 
p_5(1)(43) <= p_4(3)(43); 
p_5(1)(44) <= p_4(3)(44); 
p_5(1)(45) <= p_4(3)(45); 
p_5(1)(46) <= p_4(3)(46); 
p_5(1)(47) <= p_4(3)(47); 
p_5(1)(48) <= p_4(3)(48); 
p_5(1)(49) <= p_4(3)(49); 
p_5(1)(50) <= p_4(3)(50); 
p_5(1)(51) <= p_4(3)(51); 
p_5(1)(52) <= p_4(3)(52); 
p_5(1)(53) <= p_4(3)(53); 
p_5(1)(54) <= p_4(3)(54); 
p_5(1)(55) <= p_4(3)(55); 
p_5(1)(56) <= p_4(3)(56); 
p_5(1)(57) <= p_4(3)(57); 
p_5(1)(58) <= p_4(3)(58); 
p_5(1)(59) <= p_4(3)(59); 
p_5(1)(60) <= p_4(3)(60); 
p_5(1)(61) <= p_4(3)(61); 
p_6(0)(0) <= p_5(0)(0); 
p_6(0)(1) <= p_5(0)(1); 
ha_5_2_0: Half_Adder port map( a => p_5(0)(2), b => p_5(1)(2), cout => p_6(1)(3), s => p_6(0)(2)); 
ha_5_3_0: Half_Adder port map( a => p_5(0)(3), b => p_5(1)(3), cout => p_6(1)(4), s => p_6(0)(3)); 
fa_5_4_0: Full_Adder port map( a => p_5(0)(4), b => p_5(1)(4), cin => p_5(2)(4), cout => p_6(1)(5), s => p_6(0)(4)); 
fa_5_5_0: Full_Adder port map( a => p_5(0)(5), b => p_5(1)(5), cin => p_5(2)(5), cout => p_6(1)(6), s => p_6(0)(5)); 
fa_5_6_0: Full_Adder port map( a => p_5(0)(6), b => p_5(1)(6), cin => p_5(2)(6), cout => p_6(1)(7), s => p_6(0)(6)); 
fa_5_7_0: Full_Adder port map( a => p_5(0)(7), b => p_5(1)(7), cin => p_5(2)(7), cout => p_6(1)(8), s => p_6(0)(7)); 
fa_5_8_0: Full_Adder port map( a => p_5(0)(8), b => p_5(1)(8), cin => p_5(2)(8), cout => p_6(1)(9), s => p_6(0)(8)); 
fa_5_9_0: Full_Adder port map( a => p_5(0)(9), b => p_5(1)(9), cin => p_5(2)(9), cout => p_6(1)(10), s => p_6(0)(9)); 
fa_5_10_0: Full_Adder port map( a => p_5(0)(10), b => p_5(1)(10), cin => p_5(2)(10), cout => p_6(1)(11), s => p_6(0)(10)); 
fa_5_11_0: Full_Adder port map( a => p_5(0)(11), b => p_5(1)(11), cin => p_5(2)(11), cout => p_6(1)(12), s => p_6(0)(11)); 
fa_5_12_0: Full_Adder port map( a => p_5(0)(12), b => p_5(1)(12), cin => p_5(2)(12), cout => p_6(1)(13), s => p_6(0)(12)); 
fa_5_13_0: Full_Adder port map( a => p_5(0)(13), b => p_5(1)(13), cin => p_5(2)(13), cout => p_6(1)(14), s => p_6(0)(13)); 
fa_5_14_0: Full_Adder port map( a => p_5(0)(14), b => p_5(1)(14), cin => p_5(2)(14), cout => p_6(1)(15), s => p_6(0)(14)); 
fa_5_15_0: Full_Adder port map( a => p_5(0)(15), b => p_5(1)(15), cin => p_5(2)(15), cout => p_6(1)(16), s => p_6(0)(15)); 
fa_5_16_0: Full_Adder port map( a => p_5(0)(16), b => p_5(1)(16), cin => p_5(2)(16), cout => p_6(1)(17), s => p_6(0)(16)); 
fa_5_17_0: Full_Adder port map( a => p_5(0)(17), b => p_5(1)(17), cin => p_5(2)(17), cout => p_6(1)(18), s => p_6(0)(17)); 
fa_5_18_0: Full_Adder port map( a => p_5(0)(18), b => p_5(1)(18), cin => p_5(2)(18), cout => p_6(1)(19), s => p_6(0)(18)); 
fa_5_19_0: Full_Adder port map( a => p_5(0)(19), b => p_5(1)(19), cin => p_5(2)(19), cout => p_6(1)(20), s => p_6(0)(19)); 
fa_5_20_0: Full_Adder port map( a => p_5(0)(20), b => p_5(1)(20), cin => p_5(2)(20), cout => p_6(1)(21), s => p_6(0)(20)); 
fa_5_21_0: Full_Adder port map( a => p_5(0)(21), b => p_5(1)(21), cin => p_5(2)(21), cout => p_6(1)(22), s => p_6(0)(21)); 
fa_5_22_0: Full_Adder port map( a => p_5(0)(22), b => p_5(1)(22), cin => p_5(2)(22), cout => p_6(1)(23), s => p_6(0)(22)); 
fa_5_23_0: Full_Adder port map( a => p_5(0)(23), b => p_5(1)(23), cin => p_5(2)(23), cout => p_6(1)(24), s => p_6(0)(23)); 
fa_5_24_0: Full_Adder port map( a => p_5(0)(24), b => p_5(1)(24), cin => p_5(2)(24), cout => p_6(1)(25), s => p_6(0)(24)); 
fa_5_25_0: Full_Adder port map( a => p_5(0)(25), b => p_5(1)(25), cin => p_5(2)(25), cout => p_6(1)(26), s => p_6(0)(25)); 
fa_5_26_0: Full_Adder port map( a => p_5(0)(26), b => p_5(1)(26), cin => p_5(2)(26), cout => p_6(1)(27), s => p_6(0)(26)); 
fa_5_27_0: Full_Adder port map( a => p_5(0)(27), b => p_5(1)(27), cin => p_5(2)(27), cout => p_6(1)(28), s => p_6(0)(27)); 
fa_5_28_0: Full_Adder port map( a => p_5(0)(28), b => p_5(1)(28), cin => p_5(2)(28), cout => p_6(1)(29), s => p_6(0)(28)); 
fa_5_29_0: Full_Adder port map( a => p_5(0)(29), b => p_5(1)(29), cin => p_5(2)(29), cout => p_6(1)(30), s => p_6(0)(29)); 
fa_5_30_0: Full_Adder port map( a => p_5(0)(30), b => p_5(1)(30), cin => p_5(2)(30), cout => p_6(1)(31), s => p_6(0)(30)); 
fa_5_31_0: Full_Adder port map( a => p_5(0)(31), b => p_5(1)(31), cin => p_5(2)(31), cout => p_6(1)(32), s => p_6(0)(31)); 
fa_5_32_0: Full_Adder port map( a => p_5(0)(32), b => p_5(1)(32), cin => p_5(2)(32), cout => p_6(1)(33), s => p_6(0)(32)); 
fa_5_33_0: Full_Adder port map( a => p_5(0)(33), b => p_5(1)(33), cin => p_5(2)(33), cout => p_6(1)(34), s => p_6(0)(33)); 
fa_5_34_0: Full_Adder port map( a => p_5(0)(34), b => p_5(1)(34), cin => p_5(2)(34), cout => p_6(1)(35), s => p_6(0)(34)); 
fa_5_35_0: Full_Adder port map( a => p_5(0)(35), b => p_5(1)(35), cin => p_5(2)(35), cout => p_6(1)(36), s => p_6(0)(35)); 
fa_5_36_0: Full_Adder port map( a => p_5(0)(36), b => p_5(1)(36), cin => p_5(2)(36), cout => p_6(1)(37), s => p_6(0)(36)); 
fa_5_37_0: Full_Adder port map( a => p_5(0)(37), b => p_5(1)(37), cin => p_5(2)(37), cout => p_6(1)(38), s => p_6(0)(37)); 
fa_5_38_0: Full_Adder port map( a => p_5(0)(38), b => p_5(1)(38), cin => p_5(2)(38), cout => p_6(1)(39), s => p_6(0)(38)); 
fa_5_39_0: Full_Adder port map( a => p_5(0)(39), b => p_5(1)(39), cin => p_5(2)(39), cout => p_6(1)(40), s => p_6(0)(39)); 
fa_5_40_0: Full_Adder port map( a => p_5(0)(40), b => p_5(1)(40), cin => p_5(2)(40), cout => p_6(1)(41), s => p_6(0)(40)); 
fa_5_41_0: Full_Adder port map( a => p_5(0)(41), b => p_5(1)(41), cin => p_5(2)(41), cout => p_6(1)(42), s => p_6(0)(41)); 
fa_5_42_0: Full_Adder port map( a => p_5(0)(42), b => p_5(1)(42), cin => p_5(2)(42), cout => p_6(1)(43), s => p_6(0)(42)); 
fa_5_43_0: Full_Adder port map( a => p_5(0)(43), b => p_5(1)(43), cin => p_5(2)(43), cout => p_6(1)(44), s => p_6(0)(43)); 
fa_5_44_0: Full_Adder port map( a => p_5(0)(44), b => p_5(1)(44), cin => p_5(2)(44), cout => p_6(1)(45), s => p_6(0)(44)); 
fa_5_45_0: Full_Adder port map( a => p_5(0)(45), b => p_5(1)(45), cin => p_5(2)(45), cout => p_6(1)(46), s => p_6(0)(45)); 
fa_5_46_0: Full_Adder port map( a => p_5(0)(46), b => p_5(1)(46), cin => p_5(2)(46), cout => p_6(1)(47), s => p_6(0)(46)); 
fa_5_47_0: Full_Adder port map( a => p_5(0)(47), b => p_5(1)(47), cin => p_5(2)(47), cout => p_6(1)(48), s => p_6(0)(47)); 
fa_5_48_0: Full_Adder port map( a => p_5(0)(48), b => p_5(1)(48), cin => p_5(2)(48), cout => p_6(1)(49), s => p_6(0)(48)); 
fa_5_49_0: Full_Adder port map( a => p_5(0)(49), b => p_5(1)(49), cin => p_5(2)(49), cout => p_6(1)(50), s => p_6(0)(49)); 
fa_5_50_0: Full_Adder port map( a => p_5(0)(50), b => p_5(1)(50), cin => p_5(2)(50), cout => p_6(1)(51), s => p_6(0)(50)); 
fa_5_51_0: Full_Adder port map( a => p_5(0)(51), b => p_5(1)(51), cin => p_5(2)(51), cout => p_6(1)(52), s => p_6(0)(51)); 
fa_5_52_0: Full_Adder port map( a => p_5(0)(52), b => p_5(1)(52), cin => p_5(2)(52), cout => p_6(1)(53), s => p_6(0)(52)); 
fa_5_53_0: Full_Adder port map( a => p_5(0)(53), b => p_5(1)(53), cin => p_5(2)(53), cout => p_6(1)(54), s => p_6(0)(53)); 
fa_5_54_0: Full_Adder port map( a => p_5(0)(54), b => p_5(1)(54), cin => p_5(2)(54), cout => p_6(1)(55), s => p_6(0)(54)); 
fa_5_55_0: Full_Adder port map( a => p_5(0)(55), b => p_5(1)(55), cin => p_5(2)(55), cout => p_6(1)(56), s => p_6(0)(55)); 
fa_5_56_0: Full_Adder port map( a => p_5(0)(56), b => p_5(1)(56), cin => p_5(2)(56), cout => p_6(1)(57), s => p_6(0)(56)); 
fa_5_57_0: Full_Adder port map( a => p_5(0)(57), b => p_5(1)(57), cin => p_5(2)(57), cout => p_6(1)(58), s => p_6(0)(57)); 
fa_5_58_0: Full_Adder port map( a => p_5(0)(58), b => p_5(1)(58), cin => p_5(2)(58), cout => p_6(1)(59), s => p_6(0)(58)); 
fa_5_59_0: Full_Adder port map( a => p_5(0)(59), b => p_5(1)(59), cin => p_5(2)(59), cout => p_6(1)(60), s => p_6(0)(59)); 
fa_5_60_0: Full_Adder port map( a => p_5(0)(60), b => p_5(1)(60), cin => p_5(2)(60), cout => p_6(1)(61), s => p_6(0)(60)); 
fa_5_61_0: Full_Adder port map( a => p_5(0)(61), b => p_5(1)(61), cin => p_5(2)(61), cout => p_6(1)(62), s => p_6(0)(61)); 
fa_5_62_0: Full_Adder port map( a => p_5(0)(62), b => p_5(1)(62), cin => p_5(2)(62), cout => p_6(1)(63), s => p_6(0)(62)); 
fa_5_63_0: Full_Adder port map( a => p_5(0)(63), b => p_5(1)(63), cin => p_5(2)(63), cout => p_6(1)(64), s => p_6(0)(63)); 
p_6(1)(0) <= p_5(1)(0); 
p_6(1)(2) <= p_5(2)(2); 



END struct;
