library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
use ieee.std_logic_textio.all;

library std;
use std.textio.all;
-- entity for writing 3 samples every clock cycle
entity data_sink is
  port (
    CLK   : in std_logic;
    RST_n : in std_logic;
    VIN   : in std_logic;
	DIN_x   : in std_logic_vector(9 downto 0);
	DIN_y   : in std_logic_vector(9 downto 0);
    DIN_z   : in std_logic_vector(9 downto 0));
end data_sink;

architecture beh of data_sink is

begin  -- beh

  process (CLK, RST_n)
    file res_fp : text open WRITE_MODE is "./resultsVHDL_parallel.txt";
    variable line_out : line;    
  begin  -- process
    if RST_n = '0' then                 -- asynchronous reset (active low)
      null;
    elsif CLK'event and CLK = '1' then  -- rising clock edge
      if (VIN = '1') then
        write(line_out, conv_integer(signed(DIN_x)));
        writeline(res_fp, line_out);
		write(line_out, conv_integer(signed(DIN_y)));
        writeline(res_fp, line_out);
		write(line_out, conv_integer(signed(DIN_z)));
        writeline(res_fp, line_out);
      end if;
    end if;
  end process;

end beh;
